VERSION 5.7 ;
BUSBITCHARS "[]" ; 
DIVIDERCHAR "/" ;

UNITS
    DATABASE MICRONS 2000 ;
END UNITS

MANUFACTURINGGRID 0.007500 ;

SITE CoreSite
    SIZE 0.210 BY 1.050 ;
    CLASS CORE ;
    SYMMETRY Y ;
END CoreSite

LAYER CO
    TYPE CUT ;
END CO

LAYER M1
    TYPE ROUTING ;
    DIRECTION HORIZONTAL ;
    PITCH 0.15 0.150 ;
    OFFSET 0.000 0.000 ;
    WIDTH 0.050000 ;
END M1

LAYER VIA1
    TYPE CUT ;
END VIA1

LAYER M2
    TYPE ROUTING ;
    DIRECTION VERTICAL ;
    PITCH 0.21 0.150 ;
    OFFSET 0.105 0.000 ;
    WIDTH 0.050000 ;
END M2

LAYER VIA2
    TYPE CUT ;
END VIA2

LAYER M3
    TYPE ROUTING ;
    DIRECTION HORIZONTAL ;
    PITCH 0.150 0.150 ;
    OFFSET 0.000 0.000 ;
    WIDTH 0.050000 ;
END M3

LAYER VIA3
    TYPE CUT ;
END VIA3

LAYER M4
    TYPE ROUTING ;
    DIRECTION VERTICAL ;
    PITCH 0.150 0.150 ;
    OFFSET 0.000 0.000 ;
    WIDTH 0.050000 ;
END M4

LAYER VIA4
    TYPE CUT ;
END VIA4

LAYER M5
    TYPE ROUTING ;
    DIRECTION HORIZONTAL ;
    PITCH 0.150 0.150 ;
    OFFSET 0.000 0.000 ;
    WIDTH 0.050000 ;
END M5

LAYER VIA5
    TYPE CUT ;
END VIA5

LAYER M6
    TYPE ROUTING ;
    DIRECTION VERTICAL ;
    PITCH 0.150 0.150 ;
    OFFSET 0.000 0.000 ;
    WIDTH 0.050000 ;
END M6

LAYER VIA6
    TYPE CUT ;
END VIA6

LAYER M7
    TYPE ROUTING ;
    DIRECTION HORIZONTAL ;
    PITCH 0.120000 0.120000 ;
    OFFSET 0.000000 0.000000 ;
    WIDTH 0.600000 ;
END M7

LAYER VIA7
    TYPE CUT ;
END VIA7

LAYER M8
    TYPE ROUTING ;
    DIRECTION VERTICAL ;
    PITCH 4.5 ;
    OFFSET 0 ;
    HEIGHT 1.825 ;
    THICKNESS 3.5 ;
    FILLACTIVESPACING 3 ;
    WIDTH 3.0 ;
END M8

LAYER RV
    TYPE CUT ;
END RV

LAYER AP
    TYPE ROUTING ;
    DIRECTION HORIZONTAL ;
    PITCH   6.250000 6.250000 ;
    OFFSET 0.000000 0.000000 ;
    WIDTH   3.000000 ;

END AP

VIA VIA12_square
	RESISTANCE 12.000000 ;
	LAYER M1 ;
		RECT -0.037500 -0.037500 0.037500 0.025 ;
	LAYER VIA1 ;
		RECT -0.037500 -0.037500 0.037500 0.025 ;
	LAYER M2 ;
		RECT -0.037500 -0.037500 0.037500 0.025 ;
END VIA12_square

VIA VIA12_slot
	RESISTANCE 6.750000 ;
	LAYER M1 ;
		RECT -0.097500 -0.037500 0.097500 0.025 ;
	LAYER VIA1 ;
		RECT -0.097500 -0.037500 0.097500 0.025 ;
	LAYER M2 ;
		RECT -0.097500 -0.037500 0.097500 0.025 ;
END VIA12_slot

VIA VIA12_slotV
	RESISTANCE 6.750000 ;
	LAYER M1 ;
		RECT -0.037500 -0.097500 0.037500 0.065 ;
	LAYER VIA1 ;
		RECT -0.037500 -0.097500 0.037500 0.065 ;
	LAYER M2 ;
		RECT -0.037500 -0.097500 0.037500 0.065 ;
END VIA12_slotV

VIA VIA12_1cut DEFAULT
	RESISTANCE 12.000000 ;
	LAYER M1 ;
		RECT -0.082500 -0.037500 0.082500 0.025 ;
	LAYER VIA1 ;
		RECT -0.037500 -0.037500 0.037500 0.025 ;
	LAYER M2 ;
		RECT -0.037500 -0.082500 0.037500 0.055 ;
END VIA12_1cut

VIA VIA12_1cut_FAT_C DEFAULT
	RESISTANCE 12.000000 ;
	LAYER M1 ;
		RECT -0.112500 -0.037500 0.112500 0.025 ;
	LAYER VIA1 ;
		RECT -0.037500 -0.037500 0.037500 0.025 ;
	LAYER M2 ;
		RECT -0.037500 -0.112500 0.037500 0.075 ;
END VIA12_1cut_FAT_C

VIA VIA12_1cut_H DEFAULT
	RESISTANCE 12.000000 ;
	LAYER M1 ;
		RECT -0.082500 -0.037500 0.082500 0.025 ;
	LAYER VIA1 ;
		RECT -0.037500 -0.037500 0.037500 0.025 ;
	LAYER M2 ;
		RECT -0.082500 -0.037500 0.082500 0.025 ;
END VIA12_1cut_H

VIA VIA12_1cut_V DEFAULT
	RESISTANCE 12.000000 ;
	LAYER M1 ;
		RECT -0.037500 -0.082500 0.037500 0.055 ;
	LAYER VIA1 ;
		RECT -0.037500 -0.037500 0.037500 0.025 ;
	LAYER M2 ;
		RECT -0.037500 -0.082500 0.037500 0.055 ;
END VIA12_1cut_V

VIA VIA12_1cut_EN1415 DEFAULT
	RESISTANCE 12.000000 ;
	LAYER M1 ;
		RECT -0.075000 -0.052500 0.075000 0.035 ;
	LAYER VIA1 ;
		RECT -0.037500 -0.037500 0.037500 0.025 ;
	LAYER M2 ;
		RECT -0.052500 -0.075000 0.052500 0.05 ;
END VIA12_1cut_EN1415

VIA VIA12_2cut_P1_E DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M1 ;
		RECT -0.082500 -0.037500 0.232500 0.025 ;
	LAYER VIA1 ;
		RECT -0.022500 -0.037500 0.172500 0.025 ;
	LAYER M2 ;
		RECT -0.037500 -0.082500 0.187500 0.055 ;
END VIA12_2cut_P1_E

VIA VIA12_2cut_P1_N DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M1 ;
		RECT -0.037500 -0.082500 0.037500 0.155 ;
	LAYER VIA1 ;
		RECT -0.037500 -0.022500 0.037500 0.115 ;
	LAYER M2 ;
		RECT -0.082500 -0.037500 0.082500 0.125 ;
END VIA12_2cut_P1_N

VIA VIA12_2cut_P1_S DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M1 ;
		RECT -0.037500 -0.232500 0.037500 0.055 ;
	LAYER VIA1 ;
		RECT -0.037500 -0.172500 0.037500 0.015 ;
	LAYER M2 ;
		RECT -0.082500 -0.187500 0.082500 0.025 ;
END VIA12_2cut_P1_S

VIA VIA12_2cut_P1_W DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M1 ;
		RECT -0.232500 -0.037500 0.082500 0.025 ;
	LAYER VIA1 ;
		RECT -0.172500 -0.037500 0.022500 0.025 ;
	LAYER M2 ;
		RECT -0.187500 -0.082500 0.037500 0.055 ;
END VIA12_2cut_P1_W

VIA VIA12_2cut_P2_BLC DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M1 ;
		RECT -0.082500 -0.112500 0.082500 0.075 ;
	LAYER VIA1 ;
		RECT -0.037500 -0.097500 0.037500 0.065 ;
	LAYER M2 ;
		RECT -0.037500 -0.330000 0.037500 0.22 ;
END VIA12_2cut_P2_BLC

VIA VIA12_2cut_P2_SLN DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M1 ;
		RECT -0.082500 -0.037500 0.082500 0.125 ;
	LAYER VIA1 ;
		RECT -0.037500 -0.022500 0.037500 0.115 ;
	LAYER M2 ;
		RECT -0.037500 -0.097500 0.037500 0.375 ;
END VIA12_2cut_P2_SLN

VIA VIA12_2cut_P2_SLS DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M1 ;
		RECT -0.082500 -0.187500 0.082500 0.025 ;
	LAYER VIA1 ;
		RECT -0.037500 -0.172500 0.037500 0.015 ;
	LAYER M2 ;
		RECT -0.037500 -0.562500 0.037500 0.065 ;
END VIA12_2cut_P2_SLS

VIA VIA12_2cut_P3_CV DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M1 ;
		RECT -0.082500 -0.112500 0.082500 0.075 ;
	LAYER VIA1 ;
		RECT -0.037500 -0.097500 0.037500 0.065 ;
	LAYER M2 ;
		RECT -0.037500 -0.157500 0.037500 0.105 ;
END VIA12_2cut_P3_CV

VIA VIA12_2cut_P3_NS DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M1 ;
		RECT -0.082500 -0.037500 0.082500 0.125 ;
	LAYER VIA1 ;
		RECT -0.037500 -0.022500 0.037500 0.115 ;
	LAYER M2 ;
		RECT -0.037500 -0.082500 0.037500 0.155 ;
END VIA12_2cut_P3_NS

VIA VIA12_2cut_P3_SS DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M1 ;
		RECT -0.082500 -0.187500 0.082500 0.025 ;
	LAYER VIA1 ;
		RECT -0.037500 -0.172500 0.037500 0.015 ;
	LAYER M2 ;
		RECT -0.037500 -0.232500 0.037500 0.055 ;
END VIA12_2cut_P3_SS

VIA VIA12_4cut DEFAULT
	RESISTANCE 3.000000 ;
	LAYER M1 ;
		RECT -0.180000 -0.135000 0.180000 0.09 ;
	LAYER VIA1 ;
		RECT -0.135000 -0.135000 -0.060000 -0.04 ;
		RECT 0.060000 -0.135000 0.135000 -0.04 ;
		RECT -0.135000 0.060000 -0.060000 0.09 ;
		RECT 0.060000 0.060000 0.135000 0.09 ;
	LAYER M2 ;
		RECT -0.135000 -0.180000 0.135000 0.12 ;
END VIA12_4cut

VIA VIA12_FBD_XEN DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M1 ;
		RECT -0.037500 -0.037500 0.247500 0.085 ;
	LAYER VIA1 ;
		RECT 0.007500 0.007500 0.202500 0.055 ;
	LAYER M2 ;
		RECT -0.037500 -0.037500 0.247500 0.085 ;
END VIA12_FBD_XEN

VIA VIA12_FBD_XES DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M1 ;
		RECT -0.037500 -0.127500 0.247500 0.025 ;
	LAYER VIA1 ;
		RECT 0.007500 -0.082500 0.202500 -0.005 ;
	LAYER M2 ;
		RECT -0.037500 -0.127500 0.247500 0.025 ;
END VIA12_FBD_XES

VIA VIA12_FBD_XWN DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M1 ;
		RECT -0.247500 -0.037500 0.037500 0.085 ;
	LAYER VIA1 ;
		RECT -0.202500 0.007500 -0.007500 0.055 ;
	LAYER M2 ;
		RECT -0.247500 -0.037500 0.037500 0.085 ;
END VIA12_FBD_XWN

VIA VIA12_FBD_XWS DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M1 ;
		RECT -0.247500 -0.127500 0.037500 0.025 ;
	LAYER VIA1 ;
		RECT -0.202500 -0.082500 -0.007500 -0.005 ;
	LAYER M2 ;
		RECT -0.247500 -0.127500 0.037500 0.025 ;
END VIA12_FBD_XWS

VIA VIA12_FBD_YEN DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M1 ;
		RECT -0.037500 -0.037500 0.127500 0.165 ;
	LAYER VIA1 ;
		RECT 0.007500 0.007500 0.082500 0.135 ;
	LAYER M2 ;
		RECT -0.037500 -0.037500 0.127500 0.165 ;
END VIA12_FBD_YEN

VIA VIA12_FBD_YES DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M1 ;
		RECT -0.037500 -0.247500 0.127500 0.025 ;
	LAYER VIA1 ;
		RECT 0.007500 -0.202500 0.082500 -0.005 ;
	LAYER M2 ;
		RECT -0.037500 -0.247500 0.127500 0.025 ;
END VIA12_FBD_YES

VIA VIA12_FBD_YWN DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M1 ;
		RECT -0.127500 -0.037500 0.037500 0.165 ;
	LAYER VIA1 ;
		RECT -0.082500 0.007500 -0.007500 0.135 ;
	LAYER M2 ;
		RECT -0.127500 -0.037500 0.037500 0.165 ;
END VIA12_FBD_YWN

VIA VIA12_FBD_YWS DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M1 ;
		RECT -0.127500 -0.247500 0.037500 0.025 ;
	LAYER VIA1 ;
		RECT -0.082500 -0.202500 -0.007500 -0.005 ;
	LAYER M2 ;
		RECT -0.127500 -0.247500 0.037500 0.025 ;
END VIA12_FBD_YWS

VIA VIA12_FBS_EN DEFAULT
	RESISTANCE 12.000000 ;
	LAYER M1 ;
		RECT -0.037500 -0.037500 0.127500 0.085 ;
	LAYER VIA1 ;
		RECT 0.007500 0.007500 0.082500 0.055 ;
	LAYER M2 ;
		RECT -0.037500 -0.037500 0.127500 0.085 ;
END VIA12_FBS_EN

VIA VIA12_FBS_ES DEFAULT
	RESISTANCE 12.000000 ;
	LAYER M1 ;
		RECT -0.037500 -0.127500 0.127500 0.025 ;
	LAYER VIA1 ;
		RECT 0.007500 -0.082500 0.082500 -0.005 ;
	LAYER M2 ;
		RECT -0.037500 -0.127500 0.127500 0.025 ;
END VIA12_FBS_ES

VIA VIA12_FBS_WN DEFAULT
	RESISTANCE 12.000000 ;
	LAYER M1 ;
		RECT -0.127500 -0.037500 0.037500 0.085 ;
	LAYER VIA1 ;
		RECT -0.082500 0.007500 -0.007500 0.055 ;
	LAYER M2 ;
		RECT -0.127500 -0.037500 0.037500 0.085 ;
END VIA12_FBS_WN

VIA VIA12_FBS_WS DEFAULT
	RESISTANCE 12.000000 ;
	LAYER M1 ;
		RECT -0.127500 -0.127500 0.037500 0.025 ;
	LAYER VIA1 ;
		RECT -0.082500 -0.082500 -0.007500 -0.005 ;
	LAYER M2 ;
		RECT -0.127500 -0.127500 0.037500 0.025 ;
END VIA12_FBS_WS

VIA VIA12_PBD_E DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M1 ;
		RECT -0.052500 -0.037500 0.262500 0.025 ;
	LAYER VIA1 ;
		RECT 0.007500 -0.037500 0.202500 0.025 ;
	LAYER M2 ;
		RECT -0.037500 -0.082500 0.247500 0.055 ;
END VIA12_PBD_E

VIA VIA12_PBD_N DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M1 ;
		RECT -0.037500 -0.052500 0.037500 0.175 ;
	LAYER VIA1 ;
		RECT -0.037500 0.007500 0.037500 0.135 ;
	LAYER M2 ;
		RECT -0.082500 -0.037500 0.082500 0.165 ;
END VIA12_PBD_N

VIA VIA12_PBD_S DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M1 ;
		RECT -0.037500 -0.262500 0.037500 0.035 ;
	LAYER VIA1 ;
		RECT -0.037500 -0.202500 0.037500 -0.005 ;
	LAYER M2 ;
		RECT -0.082500 -0.247500 0.082500 0.025 ;
END VIA12_PBD_S

VIA VIA12_PBD_W DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M1 ;
		RECT -0.262500 -0.037500 0.052500 0.025 ;
	LAYER VIA1 ;
		RECT -0.202500 -0.037500 -0.007500 0.025 ;
	LAYER M2 ;
		RECT -0.247500 -0.082500 0.037500 0.055 ;
END VIA12_PBD_W

VIA VIA12_PBS_H DEFAULT
	RESISTANCE 12.000000 ;
	LAYER M1 ;
		RECT -0.082500 -0.037500 0.082500 0.025 ;
	LAYER VIA1 ;
		RECT -0.037500 -0.037500 0.037500 0.025 ;
	LAYER M2 ;
		RECT -0.082500 -0.082500 0.082500 0.055 ;
END VIA12_PBS_H

VIA VIA12_FBD20_XEN DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M1 ;
		RECT -0.037500 -0.037500 0.217500 0.065 ;
	LAYER VIA1 ;
		RECT -0.007500 -0.007500 0.187500 0.045 ;
	LAYER M2 ;
		RECT -0.037500 -0.037500 0.217500 0.065 ;
END VIA12_FBD20_XEN

VIA VIA12_FBD20_XES DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M1 ;
		RECT -0.037500 -0.097500 0.217500 0.025 ;
	LAYER VIA1 ;
		RECT -0.007500 -0.067500 0.187500 0.005 ;
	LAYER M2 ;
		RECT -0.037500 -0.097500 0.217500 0.025 ;
END VIA12_FBD20_XES

VIA VIA12_FBD20_XWN DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M1 ;
		RECT -0.217500 -0.037500 0.037500 0.065 ;
	LAYER VIA1 ;
		RECT -0.187500 -0.007500 0.007500 0.045 ;
	LAYER M2 ;
		RECT -0.217500 -0.037500 0.037500 0.065 ;
END VIA12_FBD20_XWN

VIA VIA12_FBD20_XWS DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M1 ;
		RECT -0.217500 -0.097500 0.037500 0.025 ;
	LAYER VIA1 ;
		RECT -0.187500 -0.067500 0.007500 0.005 ;
	LAYER M2 ;
		RECT -0.217500 -0.097500 0.037500 0.025 ;
END VIA12_FBD20_XWS

VIA VIA12_FBD20_YEN DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M1 ;
		RECT -0.037500 -0.037500 0.097500 0.145 ;
	LAYER VIA1 ;
		RECT -0.007500 -0.007500 0.067500 0.125 ;
	LAYER M2 ;
		RECT -0.037500 -0.037500 0.097500 0.145 ;
END VIA12_FBD20_YEN

VIA VIA12_FBD20_YES DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M1 ;
		RECT -0.037500 -0.217500 0.097500 0.025 ;
	LAYER VIA1 ;
		RECT -0.007500 -0.187500 0.067500 0.005 ;
	LAYER M2 ;
		RECT -0.037500 -0.217500 0.097500 0.025 ;
END VIA12_FBD20_YES

VIA VIA12_FBD20_YWN DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M1 ;
		RECT -0.097500 -0.037500 0.037500 0.145 ;
	LAYER VIA1 ;
		RECT -0.067500 -0.007500 0.007500 0.125 ;
	LAYER M2 ;
		RECT -0.097500 -0.037500 0.037500 0.145 ;
END VIA12_FBD20_YWN

VIA VIA12_FBD20_YWS DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M1 ;
		RECT -0.097500 -0.217500 0.037500 0.025 ;
	LAYER VIA1 ;
		RECT -0.067500 -0.187500 0.007500 0.005 ;
	LAYER M2 ;
		RECT -0.097500 -0.217500 0.037500 0.025 ;
END VIA12_FBD20_YWS

VIA VIA12_FBD30_XEN DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M1 ;
		RECT -0.037500 -0.037500 0.187500 0.085 ;
	LAYER VIA1 ;
		RECT -0.022500 0.007500 0.172500 0.055 ;
	LAYER M2 ;
		RECT -0.037500 -0.037500 0.187500 0.085 ;
END VIA12_FBD30_XEN

VIA VIA12_FBD30_XES DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M1 ;
		RECT -0.037500 -0.127500 0.187500 0.025 ;
	LAYER VIA1 ;
		RECT -0.022500 -0.082500 0.172500 -0.005 ;
	LAYER M2 ;
		RECT -0.037500 -0.127500 0.187500 0.025 ;
END VIA12_FBD30_XES

VIA VIA12_FBD30_XWN DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M1 ;
		RECT -0.187500 -0.037500 0.037500 0.085 ;
	LAYER VIA1 ;
		RECT -0.172500 0.007500 0.022500 0.055 ;
	LAYER M2 ;
		RECT -0.187500 -0.037500 0.037500 0.085 ;
END VIA12_FBD30_XWN

VIA VIA12_FBD30_XWS DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M1 ;
		RECT -0.187500 -0.127500 0.037500 0.025 ;
	LAYER VIA1 ;
		RECT -0.172500 -0.082500 0.022500 -0.005 ;
	LAYER M2 ;
		RECT -0.187500 -0.127500 0.037500 0.025 ;
END VIA12_FBD30_XWS

VIA VIA12_FBD30_YEN DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M1 ;
		RECT -0.037500 -0.037500 0.127500 0.125 ;
	LAYER VIA1 ;
		RECT 0.007500 -0.022500 0.082500 0.115 ;
	LAYER M2 ;
		RECT -0.037500 -0.037500 0.127500 0.125 ;
END VIA12_FBD30_YEN

VIA VIA12_FBD30_YES DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M1 ;
		RECT -0.037500 -0.187500 0.127500 0.025 ;
	LAYER VIA1 ;
		RECT 0.007500 -0.172500 0.082500 0.015 ;
	LAYER M2 ;
		RECT -0.037500 -0.187500 0.127500 0.025 ;
END VIA12_FBD30_YES

VIA VIA12_FBD30_YWN DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M1 ;
		RECT -0.127500 -0.037500 0.037500 0.125 ;
	LAYER VIA1 ;
		RECT -0.082500 -0.022500 -0.007500 0.115 ;
	LAYER M2 ;
		RECT -0.127500 -0.037500 0.037500 0.125 ;
END VIA12_FBD30_YWN

VIA VIA12_FBD30_YWS DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M1 ;
		RECT -0.127500 -0.187500 0.037500 0.025 ;
	LAYER VIA1 ;
		RECT -0.082500 -0.172500 -0.007500 0.015 ;
	LAYER M2 ;
		RECT -0.127500 -0.187500 0.037500 0.025 ;
END VIA12_FBD30_YWS

VIA VIA12_PBDB_E DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M1 ;
		RECT -0.007500 -0.067500 0.247500 0.045 ;
	LAYER VIA1 ;
		RECT 0.022500 -0.037500 0.217500 0.025 ;
	LAYER M2 ;
		RECT -0.037500 -0.037500 0.277500 0.025 ;
END VIA12_PBDB_E

VIA VIA12_PBDB_N DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M1 ;
		RECT -0.067500 -0.007500 0.067500 0.165 ;
	LAYER VIA1 ;
		RECT -0.037500 0.022500 0.037500 0.145 ;
	LAYER M2 ;
		RECT -0.037500 -0.037500 0.037500 0.185 ;
END VIA12_PBDB_N

VIA VIA12_PBDB_S DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M1 ;
		RECT -0.067500 -0.247500 0.067500 0.005 ;
	LAYER VIA1 ;
		RECT -0.037500 -0.217500 0.037500 -0.015 ;
	LAYER M2 ;
		RECT -0.037500 -0.277500 0.037500 0.025 ;
END VIA12_PBDB_S

VIA VIA12_PBDB_W DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M1 ;
		RECT -0.247500 -0.067500 0.007500 0.045 ;
	LAYER VIA1 ;
		RECT -0.217500 -0.037500 -0.022500 0.025 ;
	LAYER M2 ;
		RECT -0.277500 -0.037500 0.037500 0.025 ;
END VIA12_PBDB_W

VIA VIA12_PBDU_E DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M1 ;
		RECT -0.067500 -0.037500 0.247500 0.025 ;
	LAYER VIA1 ;
		RECT -0.007500 -0.037500 0.187500 0.025 ;
	LAYER M2 ;
		RECT -0.037500 -0.067500 0.217500 0.045 ;
END VIA12_PBDU_E

VIA VIA12_PBDU_N DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M1 ;
		RECT -0.037500 -0.067500 0.037500 0.165 ;
	LAYER VIA1 ;
		RECT -0.037500 -0.007500 0.037500 0.125 ;
	LAYER M2 ;
		RECT -0.067500 -0.037500 0.067500 0.145 ;
END VIA12_PBDU_N

VIA VIA12_PBDU_S DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M1 ;
		RECT -0.037500 -0.247500 0.037500 0.045 ;
	LAYER VIA1 ;
		RECT -0.037500 -0.187500 0.037500 0.005 ;
	LAYER M2 ;
		RECT -0.067500 -0.217500 0.067500 0.025 ;
END VIA12_PBDU_S

VIA VIA12_PBDU_W DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M1 ;
		RECT -0.247500 -0.037500 0.067500 0.025 ;
	LAYER VIA1 ;
		RECT -0.187500 -0.037500 0.007500 0.025 ;
	LAYER M2 ;
		RECT -0.217500 -0.067500 0.037500 0.045 ;
END VIA12_PBDU_W

VIA VIA12_PBDE_E DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M1 ;
		RECT -0.037500 -0.037500 0.277500 0.025 ;
	LAYER VIA1 ;
		RECT 0.022500 -0.037500 0.217500 0.025 ;
	LAYER M2 ;
		RECT -0.037500 -0.037500 0.277500 0.025 ;
END VIA12_PBDE_E

VIA VIA12_PBDE_N DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M1 ;
		RECT -0.037500 -0.037500 0.037500 0.185 ;
	LAYER VIA1 ;
		RECT -0.037500 0.022500 0.037500 0.145 ;
	LAYER M2 ;
		RECT -0.037500 -0.037500 0.037500 0.185 ;
END VIA12_PBDE_N

VIA VIA12_PBDE_S DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M1 ;
		RECT -0.037500 -0.277500 0.037500 0.025 ;
	LAYER VIA1 ;
		RECT -0.037500 -0.217500 0.037500 -0.015 ;
	LAYER M2 ;
		RECT -0.037500 -0.277500 0.037500 0.025 ;
END VIA12_PBDE_S

VIA VIA12_PBDE_W DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M1 ;
		RECT -0.277500 -0.037500 0.037500 0.025 ;
	LAYER VIA1 ;
		RECT -0.217500 -0.037500 -0.022500 0.025 ;
	LAYER M2 ;
		RECT -0.277500 -0.037500 0.037500 0.025 ;
END VIA12_PBDE_W

VIA VIA12_FBS25_EN DEFAULT
	RESISTANCE 12.000000 ;
	LAYER M1 ;
		RECT -0.037500 -0.037500 0.112500 0.075 ;
	LAYER VIA1 ;
		RECT 0.000000 0.000000 0.075000 0.05 ;
	LAYER M2 ;
		RECT -0.037500 -0.037500 0.112500 0.075 ;
END VIA12_FBS25_EN

VIA VIA12_FBS25_ES DEFAULT
	RESISTANCE 12.000000 ;
	LAYER M1 ;
		RECT -0.037500 -0.112500 0.112500 0.025 ;
	LAYER VIA1 ;
		RECT 0.000000 -0.075000 0.075000 0 ;
	LAYER M2 ;
		RECT -0.037500 -0.112500 0.112500 0.025 ;
END VIA12_FBS25_ES

VIA VIA12_FBS25_WN DEFAULT
	RESISTANCE 12.000000 ;
	LAYER M1 ;
		RECT -0.112500 -0.037500 0.037500 0.075 ;
	LAYER VIA1 ;
		RECT -0.075000 0.000000 0.000000 0.05 ;
	LAYER M2 ;
		RECT -0.112500 -0.037500 0.037500 0.075 ;
END VIA12_FBS25_WN

VIA VIA12_FBS25_WS DEFAULT
	RESISTANCE 12.000000 ;
	LAYER M1 ;
		RECT -0.112500 -0.112500 0.037500 0.025 ;
	LAYER VIA1 ;
		RECT -0.075000 -0.075000 0.000000 0 ;
	LAYER M2 ;
		RECT -0.112500 -0.112500 0.037500 0.025 ;
END VIA12_FBS25_WS

VIA VIA12_PBSU_H DEFAULT
	RESISTANCE 12.000000 ;
	LAYER M1 ;
		RECT -0.082500 -0.037500 0.082500 0.025 ;
	LAYER VIA1 ;
		RECT -0.037500 -0.037500 0.037500 0.025 ;
	LAYER M2 ;
		RECT -0.052500 -0.075000 0.052500 0.05 ;
END VIA12_PBSU_H

VIA VIA12_PBSB_H DEFAULT
	RESISTANCE 12.000000 ;
	LAYER M1 ;
		RECT -0.075000 -0.052500 0.075000 0.035 ;
	LAYER VIA1 ;
		RECT -0.037500 -0.037500 0.037500 0.025 ;
	LAYER M2 ;
		RECT -0.037500 -0.082500 0.037500 0.055 ;
END VIA12_PBSB_H


VIA VIA23_1cut DEFAULT
	RESISTANCE 12.000000 ;
	LAYER M2 ;
		RECT -0.037500 -0.082500 0.037500 0.055 ;
	LAYER VIA2 ;
		RECT -0.037500 -0.037500 0.037500 0.025 ;
	LAYER M3 ;
		RECT -0.082500 -0.037500 0.082500 0.025 ;
END VIA23_1cut

VIA VIA23_1cut_FAT_C DEFAULT
	RESISTANCE 12.000000 ;
	LAYER M2 ;
		RECT -0.037500 -0.112500 0.037500 0.075 ;
	LAYER VIA2 ;
		RECT -0.037500 -0.037500 0.037500 0.025 ;
	LAYER M3 ;
		RECT -0.112500 -0.037500 0.112500 0.025 ;
END VIA23_1cut_FAT_C

VIA VIA23_1cut_EN1415 DEFAULT
	RESISTANCE 12.000000 ;
	LAYER M2 ;
		RECT -0.052500 -0.075000 0.052500 0.05 ;
	LAYER VIA2 ;
		RECT -0.037500 -0.037500 0.037500 0.025 ;
	LAYER M3 ;
		RECT -0.075000 -0.052500 0.075000 0.035 ;
END VIA23_1cut_EN1415

VIA VIA23_1stack_C DEFAULT
	RESISTANCE 12.000000 ;
	LAYER M2 ;
		RECT -0.037500 -0.210000 0.037500 0.14 ;
	LAYER VIA2 ;
		RECT -0.037500 -0.037500 0.037500 0.025 ;
	LAYER M3 ;
		RECT -0.082500 -0.037500 0.082500 0.025 ;
END VIA23_1stack_C

VIA VIA23_1stack_N DEFAULT
	RESISTANCE 12.000000 ;
	LAYER M2 ;
		RECT -0.037500 -0.082500 0.037500 0.225 ;
	LAYER VIA2 ;
		RECT -0.037500 -0.037500 0.037500 0.025 ;
	LAYER M3 ;
		RECT -0.082500 -0.037500 0.082500 0.025 ;
END VIA23_1stack_N

VIA VIA23_1stack_S DEFAULT
	RESISTANCE 12.000000 ;
	LAYER M2 ;
		RECT -0.037500 -0.337500 0.037500 0.055 ;
	LAYER VIA2 ;
		RECT -0.037500 -0.037500 0.037500 0.025 ;
	LAYER M3 ;
		RECT -0.082500 -0.037500 0.082500 0.025 ;
END VIA23_1stack_S

VIA VIA23_2cut_P1_N DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M2 ;
		RECT -0.037500 -0.082500 0.037500 0.155 ;
	LAYER VIA2 ;
		RECT -0.037500 -0.022500 0.037500 0.115 ;
	LAYER M3 ;
		RECT -0.082500 -0.037500 0.082500 0.125 ;
END VIA23_2cut_P1_N

VIA VIA23_2cut_P1_S DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M2 ;
		RECT -0.037500 -0.232500 0.037500 0.055 ;
	LAYER VIA2 ;
		RECT -0.037500 -0.172500 0.037500 0.015 ;
	LAYER M3 ;
		RECT -0.082500 -0.187500 0.082500 0.025 ;
END VIA23_2cut_P1_S

VIA VIA23_2cut_P2_BLC DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M2 ;
		RECT -0.112500 -0.082500 0.112500 0.055 ;
	LAYER VIA2 ;
		RECT -0.097500 -0.037500 0.097500 0.025 ;
	LAYER M3 ;
		RECT -0.330000 -0.037500 0.330000 0.025 ;
END VIA23_2cut_P2_BLC

VIA VIA23_2cut_P2_BLE DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M2 ;
		RECT -0.037500 -0.082500 0.187500 0.055 ;
	LAYER VIA2 ;
		RECT -0.022500 -0.037500 0.172500 0.025 ;
	LAYER M3 ;
		RECT -0.255000 -0.037500 0.405000 0.025 ;
END VIA23_2cut_P2_BLE

VIA VIA23_2cut_P2_BLW DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M2 ;
		RECT -0.187500 -0.082500 0.037500 0.055 ;
	LAYER VIA2 ;
		RECT -0.172500 -0.037500 0.022500 0.025 ;
	LAYER M3 ;
		RECT -0.405000 -0.037500 0.255000 0.025 ;
END VIA23_2cut_P2_BLW

VIA VIA23_2cut_P2_SLE DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M2 ;
		RECT -0.037500 -0.082500 0.187500 0.055 ;
	LAYER VIA2 ;
		RECT -0.022500 -0.037500 0.172500 0.025 ;
	LAYER M3 ;
		RECT -0.097500 -0.037500 0.562500 0.025 ;
END VIA23_2cut_P2_SLE

VIA VIA23_2cut_P2_SLW DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M2 ;
		RECT -0.187500 -0.082500 0.037500 0.055 ;
	LAYER VIA2 ;
		RECT -0.172500 -0.037500 0.022500 0.025 ;
	LAYER M3 ;
		RECT -0.562500 -0.037500 0.097500 0.025 ;
END VIA23_2cut_P2_SLW

VIA VIA23_2cut_P3_E DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M2 ;
		RECT -0.037500 -0.082500 0.187500 0.055 ;
	LAYER VIA2 ;
		RECT -0.022500 -0.037500 0.172500 0.025 ;
	LAYER M3 ;
		RECT -0.082500 -0.037500 0.232500 0.025 ;
END VIA23_2cut_P3_E

VIA VIA23_2cut_P3_W DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M2 ;
		RECT -0.187500 -0.082500 0.037500 0.055 ;
	LAYER VIA2 ;
		RECT -0.172500 -0.037500 0.022500 0.025 ;
	LAYER M3 ;
		RECT -0.232500 -0.037500 0.082500 0.025 ;
END VIA23_2cut_P3_W

VIA VIA23_4cut DEFAULT
	RESISTANCE 3.000000 ;
	LAYER M2 ;
		RECT -0.135000 -0.180000 0.135000 0.12 ;
	LAYER VIA2 ;
		RECT -0.135000 -0.135000 -0.060000 -0.04 ;
		RECT 0.060000 -0.135000 0.135000 -0.04 ;
		RECT -0.135000 0.060000 -0.060000 0.09 ;
		RECT 0.060000 0.060000 0.135000 0.09 ;
	LAYER M3 ;
		RECT -0.180000 -0.135000 0.180000 0.09 ;
END VIA23_4cut

VIA VIA23_FBD_XEN DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M2 ;
		RECT -0.037500 -0.037500 0.247500 0.085 ;
	LAYER VIA2 ;
		RECT 0.007500 0.007500 0.202500 0.055 ;
	LAYER M3 ;
		RECT -0.037500 -0.037500 0.247500 0.085 ;
END VIA23_FBD_XEN

VIA VIA23_FBD_XES DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M2 ;
		RECT -0.037500 -0.127500 0.247500 0.025 ;
	LAYER VIA2 ;
		RECT 0.007500 -0.082500 0.202500 -0.005 ;
	LAYER M3 ;
		RECT -0.037500 -0.127500 0.247500 0.025 ;
END VIA23_FBD_XES

VIA VIA23_FBD_XWN DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M2 ;
		RECT -0.247500 -0.037500 0.037500 0.085 ;
	LAYER VIA2 ;
		RECT -0.202500 0.007500 -0.007500 0.055 ;
	LAYER M3 ;
		RECT -0.247500 -0.037500 0.037500 0.085 ;
END VIA23_FBD_XWN

VIA VIA23_FBD_XWS DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M2 ;
		RECT -0.247500 -0.127500 0.037500 0.025 ;
	LAYER VIA2 ;
		RECT -0.202500 -0.082500 -0.007500 -0.005 ;
	LAYER M3 ;
		RECT -0.247500 -0.127500 0.037500 0.025 ;
END VIA23_FBD_XWS

VIA VIA23_FBD_YEN DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M2 ;
		RECT -0.037500 -0.037500 0.127500 0.165 ;
	LAYER VIA2 ;
		RECT 0.007500 0.007500 0.082500 0.135 ;
	LAYER M3 ;
		RECT -0.037500 -0.037500 0.127500 0.165 ;
END VIA23_FBD_YEN

VIA VIA23_FBD_YES DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M2 ;
		RECT -0.037500 -0.247500 0.127500 0.025 ;
	LAYER VIA2 ;
		RECT 0.007500 -0.202500 0.082500 -0.005 ;
	LAYER M3 ;
		RECT -0.037500 -0.247500 0.127500 0.025 ;
END VIA23_FBD_YES

VIA VIA23_FBD_YWN DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M2 ;
		RECT -0.127500 -0.037500 0.037500 0.165 ;
	LAYER VIA2 ;
		RECT -0.082500 0.007500 -0.007500 0.135 ;
	LAYER M3 ;
		RECT -0.127500 -0.037500 0.037500 0.165 ;
END VIA23_FBD_YWN

VIA VIA23_FBD_YWS DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M2 ;
		RECT -0.127500 -0.247500 0.037500 0.025 ;
	LAYER VIA2 ;
		RECT -0.082500 -0.202500 -0.007500 -0.005 ;
	LAYER M3 ;
		RECT -0.127500 -0.247500 0.037500 0.025 ;
END VIA23_FBD_YWS

VIA VIA23_FBS DEFAULT
	RESISTANCE 12.000000 ;
	LAYER M2 ;
		RECT -0.082500 -0.082500 0.082500 0.055 ;
	LAYER VIA2 ;
		RECT -0.037500 -0.037500 0.037500 0.025 ;
	LAYER M3 ;
		RECT -0.082500 -0.082500 0.082500 0.055 ;
END VIA23_FBS

VIA VIA23_FBS_EN DEFAULT
	RESISTANCE 12.000000 ;
	LAYER M2 ;
		RECT -0.037500 -0.037500 0.127500 0.085 ;
	LAYER VIA2 ;
		RECT 0.007500 0.007500 0.082500 0.055 ;
	LAYER M3 ;
		RECT -0.037500 -0.037500 0.127500 0.085 ;
END VIA23_FBS_EN

VIA VIA23_FBS_ES DEFAULT
	RESISTANCE 12.000000 ;
	LAYER M2 ;
		RECT -0.037500 -0.127500 0.127500 0.025 ;
	LAYER VIA2 ;
		RECT 0.007500 -0.082500 0.082500 -0.005 ;
	LAYER M3 ;
		RECT -0.037500 -0.127500 0.127500 0.025 ;
END VIA23_FBS_ES

VIA VIA23_FBS_WN DEFAULT
	RESISTANCE 12.000000 ;
	LAYER M2 ;
		RECT -0.127500 -0.037500 0.037500 0.085 ;
	LAYER VIA2 ;
		RECT -0.082500 0.007500 -0.007500 0.055 ;
	LAYER M3 ;
		RECT -0.127500 -0.037500 0.037500 0.085 ;
END VIA23_FBS_WN

VIA VIA23_FBS_WS DEFAULT
	RESISTANCE 12.000000 ;
	LAYER M2 ;
		RECT -0.127500 -0.127500 0.037500 0.025 ;
	LAYER VIA2 ;
		RECT -0.082500 -0.082500 -0.007500 -0.005 ;
	LAYER M3 ;
		RECT -0.127500 -0.127500 0.037500 0.025 ;
END VIA23_FBS_WS

VIA VIA23_PBD_E DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M2 ;
		RECT -0.052500 -0.037500 0.262500 0.025 ;
	LAYER VIA2 ;
		RECT 0.007500 -0.037500 0.202500 0.025 ;
	LAYER M3 ;
		RECT -0.037500 -0.082500 0.247500 0.055 ;
END VIA23_PBD_E

VIA VIA23_PBD_N DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M2 ;
		RECT -0.037500 -0.052500 0.037500 0.175 ;
	LAYER VIA2 ;
		RECT -0.037500 0.007500 0.037500 0.135 ;
	LAYER M3 ;
		RECT -0.082500 -0.037500 0.082500 0.165 ;
END VIA23_PBD_N

VIA VIA23_PBD_S DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M2 ;
		RECT -0.037500 -0.262500 0.037500 0.035 ;
	LAYER VIA2 ;
		RECT -0.037500 -0.202500 0.037500 -0.005 ;
	LAYER M3 ;
		RECT -0.082500 -0.247500 0.082500 0.025 ;
END VIA23_PBD_S

VIA VIA23_PBD_W DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M2 ;
		RECT -0.262500 -0.037500 0.052500 0.025 ;
	LAYER VIA2 ;
		RECT -0.202500 -0.037500 -0.007500 0.025 ;
	LAYER M3 ;
		RECT -0.247500 -0.082500 0.037500 0.055 ;
END VIA23_PBD_W

VIA VIA23_PBS_H DEFAULT
	RESISTANCE 12.000000 ;
	LAYER M2 ;
		RECT -0.082500 -0.037500 0.082500 0.025 ;
	LAYER VIA2 ;
		RECT -0.037500 -0.037500 0.037500 0.025 ;
	LAYER M3 ;
		RECT -0.082500 -0.082500 0.082500 0.055 ;
END VIA23_PBS_H

VIA VIA23_PBS_V DEFAULT
	RESISTANCE 12.000000 ;
	LAYER M2 ;
		RECT -0.037500 -0.082500 0.037500 0.055 ;
	LAYER VIA2 ;
		RECT -0.037500 -0.037500 0.037500 0.025 ;
	LAYER M3 ;
		RECT -0.082500 -0.082500 0.082500 0.055 ;
END VIA23_PBS_V

VIA VIA23_FBD20_XEN DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M2 ;
		RECT -0.037500 -0.037500 0.217500 0.065 ;
	LAYER VIA2 ;
		RECT -0.007500 -0.007500 0.187500 0.045 ;
	LAYER M3 ;
		RECT -0.037500 -0.037500 0.217500 0.065 ;
END VIA23_FBD20_XEN

VIA VIA23_FBD20_XES DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M2 ;
		RECT -0.037500 -0.097500 0.217500 0.025 ;
	LAYER VIA2 ;
		RECT -0.007500 -0.067500 0.187500 0.005 ;
	LAYER M3 ;
		RECT -0.037500 -0.097500 0.217500 0.025 ;
END VIA23_FBD20_XES

VIA VIA23_FBD20_XWN DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M2 ;
		RECT -0.217500 -0.037500 0.037500 0.065 ;
	LAYER VIA2 ;
		RECT -0.187500 -0.007500 0.007500 0.045 ;
	LAYER M3 ;
		RECT -0.217500 -0.037500 0.037500 0.065 ;
END VIA23_FBD20_XWN

VIA VIA23_FBD20_XWS DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M2 ;
		RECT -0.217500 -0.097500 0.037500 0.025 ;
	LAYER VIA2 ;
		RECT -0.187500 -0.067500 0.007500 0.005 ;
	LAYER M3 ;
		RECT -0.217500 -0.097500 0.037500 0.025 ;
END VIA23_FBD20_XWS

VIA VIA23_FBD20_YEN DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M2 ;
		RECT -0.037500 -0.037500 0.097500 0.145 ;
	LAYER VIA2 ;
		RECT -0.007500 -0.007500 0.067500 0.125 ;
	LAYER M3 ;
		RECT -0.037500 -0.037500 0.097500 0.145 ;
END VIA23_FBD20_YEN

VIA VIA23_FBD20_YES DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M2 ;
		RECT -0.037500 -0.217500 0.097500 0.025 ;
	LAYER VIA2 ;
		RECT -0.007500 -0.187500 0.067500 0.005 ;
	LAYER M3 ;
		RECT -0.037500 -0.217500 0.097500 0.025 ;
END VIA23_FBD20_YES

VIA VIA23_FBD20_YWN DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M2 ;
		RECT -0.097500 -0.037500 0.037500 0.145 ;
	LAYER VIA2 ;
		RECT -0.067500 -0.007500 0.007500 0.125 ;
	LAYER M3 ;
		RECT -0.097500 -0.037500 0.037500 0.145 ;
END VIA23_FBD20_YWN

VIA VIA23_FBD20_YWS DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M2 ;
		RECT -0.097500 -0.217500 0.037500 0.025 ;
	LAYER VIA2 ;
		RECT -0.067500 -0.187500 0.007500 0.005 ;
	LAYER M3 ;
		RECT -0.097500 -0.217500 0.037500 0.025 ;
END VIA23_FBD20_YWS

VIA VIA23_FBD30_XEN DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M2 ;
		RECT -0.037500 -0.037500 0.187500 0.085 ;
	LAYER VIA2 ;
		RECT -0.022500 0.007500 0.172500 0.055 ;
	LAYER M3 ;
		RECT -0.037500 -0.037500 0.187500 0.085 ;
END VIA23_FBD30_XEN

VIA VIA23_FBD30_XES DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M2 ;
		RECT -0.037500 -0.127500 0.187500 0.025 ;
	LAYER VIA2 ;
		RECT -0.022500 -0.082500 0.172500 -0.005 ;
	LAYER M3 ;
		RECT -0.037500 -0.127500 0.187500 0.025 ;
END VIA23_FBD30_XES

VIA VIA23_FBD30_XWN DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M2 ;
		RECT -0.187500 -0.037500 0.037500 0.085 ;
	LAYER VIA2 ;
		RECT -0.172500 0.007500 0.022500 0.055 ;
	LAYER M3 ;
		RECT -0.187500 -0.037500 0.037500 0.085 ;
END VIA23_FBD30_XWN

VIA VIA23_FBD30_XWS DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M2 ;
		RECT -0.187500 -0.127500 0.037500 0.025 ;
	LAYER VIA2 ;
		RECT -0.172500 -0.082500 0.022500 -0.005 ;
	LAYER M3 ;
		RECT -0.187500 -0.127500 0.037500 0.025 ;
END VIA23_FBD30_XWS

VIA VIA23_FBD30_YEN DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M2 ;
		RECT -0.037500 -0.037500 0.127500 0.125 ;
	LAYER VIA2 ;
		RECT 0.007500 -0.022500 0.082500 0.115 ;
	LAYER M3 ;
		RECT -0.037500 -0.037500 0.127500 0.125 ;
END VIA23_FBD30_YEN

VIA VIA23_FBD30_YES DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M2 ;
		RECT -0.037500 -0.187500 0.127500 0.025 ;
	LAYER VIA2 ;
		RECT 0.007500 -0.172500 0.082500 0.015 ;
	LAYER M3 ;
		RECT -0.037500 -0.187500 0.127500 0.025 ;
END VIA23_FBD30_YES

VIA VIA23_FBD30_YWN DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M2 ;
		RECT -0.127500 -0.037500 0.037500 0.125 ;
	LAYER VIA2 ;
		RECT -0.082500 -0.022500 -0.007500 0.115 ;
	LAYER M3 ;
		RECT -0.127500 -0.037500 0.037500 0.125 ;
END VIA23_FBD30_YWN

VIA VIA23_FBD30_YWS DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M2 ;
		RECT -0.127500 -0.187500 0.037500 0.025 ;
	LAYER VIA2 ;
		RECT -0.082500 -0.172500 -0.007500 0.015 ;
	LAYER M3 ;
		RECT -0.127500 -0.187500 0.037500 0.025 ;
END VIA23_FBD30_YWS

VIA VIA23_PBDB_E DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M2 ;
		RECT -0.007500 -0.067500 0.247500 0.045 ;
	LAYER VIA2 ;
		RECT 0.022500 -0.037500 0.217500 0.025 ;
	LAYER M3 ;
		RECT -0.037500 -0.037500 0.277500 0.025 ;
END VIA23_PBDB_E

VIA VIA23_PBDB_N DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M2 ;
		RECT -0.067500 -0.007500 0.067500 0.165 ;
	LAYER VIA2 ;
		RECT -0.037500 0.022500 0.037500 0.145 ;
	LAYER M3 ;
		RECT -0.037500 -0.037500 0.037500 0.185 ;
END VIA23_PBDB_N

VIA VIA23_PBDB_S DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M2 ;
		RECT -0.067500 -0.247500 0.067500 0.005 ;
	LAYER VIA2 ;
		RECT -0.037500 -0.217500 0.037500 -0.015 ;
	LAYER M3 ;
		RECT -0.037500 -0.277500 0.037500 0.025 ;
END VIA23_PBDB_S

VIA VIA23_PBDB_W DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M2 ;
		RECT -0.247500 -0.067500 0.007500 0.045 ;
	LAYER VIA2 ;
		RECT -0.217500 -0.037500 -0.022500 0.025 ;
	LAYER M3 ;
		RECT -0.277500 -0.037500 0.037500 0.025 ;
END VIA23_PBDB_W

VIA VIA23_PBDU_E DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M2 ;
		RECT -0.067500 -0.037500 0.247500 0.025 ;
	LAYER VIA2 ;
		RECT -0.007500 -0.037500 0.187500 0.025 ;
	LAYER M3 ;
		RECT -0.037500 -0.067500 0.217500 0.045 ;
END VIA23_PBDU_E

VIA VIA23_PBDU_N DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M2 ;
		RECT -0.037500 -0.067500 0.037500 0.165 ;
	LAYER VIA2 ;
		RECT -0.037500 -0.007500 0.037500 0.125 ;
	LAYER M3 ;
		RECT -0.067500 -0.037500 0.067500 0.145 ;
END VIA23_PBDU_N

VIA VIA23_PBDU_S DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M2 ;
		RECT -0.037500 -0.247500 0.037500 0.045 ;
	LAYER VIA2 ;
		RECT -0.037500 -0.187500 0.037500 0.005 ;
	LAYER M3 ;
		RECT -0.067500 -0.217500 0.067500 0.025 ;
END VIA23_PBDU_S

VIA VIA23_PBDU_W DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M2 ;
		RECT -0.247500 -0.037500 0.067500 0.025 ;
	LAYER VIA2 ;
		RECT -0.187500 -0.037500 0.007500 0.025 ;
	LAYER M3 ;
		RECT -0.217500 -0.067500 0.037500 0.045 ;
END VIA23_PBDU_W

VIA VIA23_PBDE_E DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M2 ;
		RECT -0.037500 -0.037500 0.277500 0.025 ;
	LAYER VIA2 ;
		RECT 0.022500 -0.037500 0.217500 0.025 ;
	LAYER M3 ;
		RECT -0.037500 -0.037500 0.277500 0.025 ;
END VIA23_PBDE_E

VIA VIA23_PBDE_N DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M2 ;
		RECT -0.037500 -0.037500 0.037500 0.185 ;
	LAYER VIA2 ;
		RECT -0.037500 0.022500 0.037500 0.145 ;
	LAYER M3 ;
		RECT -0.037500 -0.037500 0.037500 0.185 ;
END VIA23_PBDE_N

VIA VIA23_PBDE_S DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M2 ;
		RECT -0.037500 -0.277500 0.037500 0.025 ;
	LAYER VIA2 ;
		RECT -0.037500 -0.217500 0.037500 -0.015 ;
	LAYER M3 ;
		RECT -0.037500 -0.277500 0.037500 0.025 ;
END VIA23_PBDE_S

VIA VIA23_PBDE_W DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M2 ;
		RECT -0.277500 -0.037500 0.037500 0.025 ;
	LAYER VIA2 ;
		RECT -0.217500 -0.037500 -0.022500 0.025 ;
	LAYER M3 ;
		RECT -0.277500 -0.037500 0.037500 0.025 ;
END VIA23_PBDE_W

VIA VIA23_FBS25 DEFAULT
	RESISTANCE 12.000000 ;
	LAYER M2 ;
		RECT -0.075000 -0.075000 0.075000 0.05 ;
	LAYER VIA2 ;
		RECT -0.037500 -0.037500 0.037500 0.025 ;
	LAYER M3 ;
		RECT -0.075000 -0.075000 0.075000 0.05 ;
END VIA23_FBS25

VIA VIA23_FBS25_EN DEFAULT
	RESISTANCE 12.000000 ;
	LAYER M2 ;
		RECT -0.037500 -0.037500 0.112500 0.075 ;
	LAYER VIA2 ;
		RECT 0.000000 0.000000 0.075000 0.05 ;
	LAYER M3 ;
		RECT -0.037500 -0.037500 0.112500 0.075 ;
END VIA23_FBS25_EN

VIA VIA23_FBS25_ES DEFAULT
	RESISTANCE 12.000000 ;
	LAYER M2 ;
		RECT -0.037500 -0.112500 0.112500 0.025 ;
	LAYER VIA2 ;
		RECT 0.000000 -0.075000 0.075000 0 ;
	LAYER M3 ;
		RECT -0.037500 -0.112500 0.112500 0.025 ;
END VIA23_FBS25_ES

VIA VIA23_FBS25_WN DEFAULT
	RESISTANCE 12.000000 ;
	LAYER M2 ;
		RECT -0.112500 -0.037500 0.037500 0.075 ;
	LAYER VIA2 ;
		RECT -0.075000 0.000000 0.000000 0.05 ;
	LAYER M3 ;
		RECT -0.112500 -0.037500 0.037500 0.075 ;
END VIA23_FBS25_WN

VIA VIA23_FBS25_WS DEFAULT
	RESISTANCE 12.000000 ;
	LAYER M2 ;
		RECT -0.112500 -0.112500 0.037500 0.025 ;
	LAYER VIA2 ;
		RECT -0.075000 -0.075000 0.000000 0 ;
	LAYER M3 ;
		RECT -0.112500 -0.112500 0.037500 0.025 ;
END VIA23_FBS25_WS

VIA VIA23_PBSU_H DEFAULT
	RESISTANCE 12.000000 ;
	LAYER M2 ;
		RECT -0.082500 -0.037500 0.082500 0.025 ;
	LAYER VIA2 ;
		RECT -0.037500 -0.037500 0.037500 0.025 ;
	LAYER M3 ;
		RECT -0.052500 -0.075000 0.052500 0.05 ;
END VIA23_PBSU_H

VIA VIA23_PBSU_V DEFAULT
	RESISTANCE 12.000000 ;
	LAYER M2 ;
		RECT -0.037500 -0.082500 0.037500 0.055 ;
	LAYER VIA2 ;
		RECT -0.037500 -0.037500 0.037500 0.025 ;
	LAYER M3 ;
		RECT -0.075000 -0.052500 0.075000 0.035 ;
END VIA23_PBSU_V

VIA VIA23_PBSB_H DEFAULT
	RESISTANCE 12.000000 ;
	LAYER M2 ;
		RECT -0.075000 -0.052500 0.075000 0.035 ;
	LAYER VIA2 ;
		RECT -0.037500 -0.037500 0.037500 0.025 ;
	LAYER M3 ;
		RECT -0.037500 -0.082500 0.037500 0.055 ;
END VIA23_PBSB_H

VIA VIA23_PBSB_V DEFAULT
	RESISTANCE 12.000000 ;
	LAYER M2 ;
		RECT -0.052500 -0.075000 0.052500 0.05 ;
	LAYER VIA2 ;
		RECT -0.037500 -0.037500 0.037500 0.025 ;
	LAYER M3 ;
		RECT -0.082500 -0.037500 0.082500 0.025 ;
END VIA23_PBSB_V


VIA VIA34_1cut DEFAULT
	RESISTANCE 12.000000 ;
	LAYER M3 ;
		RECT -0.082500 -0.037500 0.082500 0.025 ;
	LAYER VIA3 ;
		RECT -0.037500 -0.037500 0.037500 0.025 ;
	LAYER M4 ;
		RECT -0.037500 -0.082500 0.037500 0.055 ;
END VIA34_1cut

VIA VIA34_1cut_FAT_C DEFAULT
	RESISTANCE 12.000000 ;
	LAYER M3 ;
		RECT -0.112500 -0.037500 0.112500 0.025 ;
	LAYER VIA3 ;
		RECT -0.037500 -0.037500 0.037500 0.025 ;
	LAYER M4 ;
		RECT -0.037500 -0.112500 0.037500 0.075 ;
END VIA34_1cut_FAT_C

VIA VIA34_1cut_EN1415 DEFAULT
	RESISTANCE 12.000000 ;
	LAYER M3 ;
		RECT -0.075000 -0.052500 0.075000 0.035 ;
	LAYER VIA3 ;
		RECT -0.037500 -0.037500 0.037500 0.025 ;
	LAYER M4 ;
		RECT -0.052500 -0.075000 0.052500 0.05 ;
END VIA34_1cut_EN1415

VIA VIA34_1stack_C DEFAULT
	RESISTANCE 12.000000 ;
	LAYER M3 ;
		RECT -0.255000 -0.037500 0.255000 0.025 ;
	LAYER VIA3 ;
		RECT -0.037500 -0.037500 0.037500 0.025 ;
	LAYER M4 ;
		RECT -0.037500 -0.082500 0.037500 0.055 ;
END VIA34_1stack_C

VIA VIA34_1stack_E DEFAULT
	RESISTANCE 12.000000 ;
	LAYER M3 ;
		RECT -0.082500 -0.037500 0.427500 0.025 ;
	LAYER VIA3 ;
		RECT -0.037500 -0.037500 0.037500 0.025 ;
	LAYER M4 ;
		RECT -0.037500 -0.082500 0.037500 0.055 ;
END VIA34_1stack_E

VIA VIA34_1stack_W DEFAULT
	RESISTANCE 12.000000 ;
	LAYER M3 ;
		RECT -0.427500 -0.037500 0.082500 0.025 ;
	LAYER VIA3 ;
		RECT -0.037500 -0.037500 0.037500 0.025 ;
	LAYER M4 ;
		RECT -0.037500 -0.082500 0.037500 0.055 ;
END VIA34_1stack_W

VIA VIA34_2cut_P1_E DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M3 ;
		RECT -0.082500 -0.037500 0.232500 0.025 ;
	LAYER VIA3 ;
		RECT -0.022500 -0.037500 0.172500 0.025 ;
	LAYER M4 ;
		RECT -0.037500 -0.082500 0.187500 0.055 ;
END VIA34_2cut_P1_E

VIA VIA34_2cut_P1_W DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M3 ;
		RECT -0.232500 -0.037500 0.082500 0.025 ;
	LAYER VIA3 ;
		RECT -0.172500 -0.037500 0.022500 0.025 ;
	LAYER M4 ;
		RECT -0.187500 -0.082500 0.037500 0.055 ;
END VIA34_2cut_P1_W

VIA VIA34_2cut_P2_BLC DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M3 ;
		RECT -0.082500 -0.112500 0.082500 0.075 ;
	LAYER VIA3 ;
		RECT -0.037500 -0.097500 0.037500 0.065 ;
	LAYER M4 ;
		RECT -0.037500 -0.330000 0.037500 0.22 ;
END VIA34_2cut_P2_BLC

VIA VIA34_2cut_P2_BLN DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M3 ;
		RECT -0.082500 -0.037500 0.082500 0.125 ;
	LAYER VIA3 ;
		RECT -0.037500 -0.022500 0.037500 0.115 ;
	LAYER M4 ;
		RECT -0.037500 -0.255000 0.037500 0.27 ;
END VIA34_2cut_P2_BLN

VIA VIA34_2cut_P2_BLS DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M3 ;
		RECT -0.082500 -0.187500 0.082500 0.025 ;
	LAYER VIA3 ;
		RECT -0.037500 -0.172500 0.037500 0.015 ;
	LAYER M4 ;
		RECT -0.037500 -0.405000 0.037500 0.17 ;
END VIA34_2cut_P2_BLS

VIA VIA34_2cut_P2_SLN DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M3 ;
		RECT -0.082500 -0.037500 0.082500 0.125 ;
	LAYER VIA3 ;
		RECT -0.037500 -0.022500 0.037500 0.115 ;
	LAYER M4 ;
		RECT -0.037500 -0.097500 0.037500 0.375 ;
END VIA34_2cut_P2_SLN

VIA VIA34_2cut_P2_SLS DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M3 ;
		RECT -0.082500 -0.187500 0.082500 0.025 ;
	LAYER VIA3 ;
		RECT -0.037500 -0.172500 0.037500 0.015 ;
	LAYER M4 ;
		RECT -0.037500 -0.562500 0.037500 0.065 ;
END VIA34_2cut_P2_SLS

VIA VIA34_2cut_P3_N DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M3 ;
		RECT -0.082500 -0.037500 0.082500 0.125 ;
	LAYER VIA3 ;
		RECT -0.037500 -0.022500 0.037500 0.115 ;
	LAYER M4 ;
		RECT -0.037500 -0.082500 0.037500 0.155 ;
END VIA34_2cut_P3_N

VIA VIA34_2cut_P3_S DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M3 ;
		RECT -0.082500 -0.187500 0.082500 0.025 ;
	LAYER VIA3 ;
		RECT -0.037500 -0.172500 0.037500 0.015 ;
	LAYER M4 ;
		RECT -0.037500 -0.232500 0.037500 0.055 ;
END VIA34_2cut_P3_S

VIA VIA34_4cut DEFAULT
	RESISTANCE 3.000000 ;
	LAYER M3 ;
		RECT -0.180000 -0.135000 0.180000 0.09 ;
	LAYER VIA3 ;
		RECT -0.135000 -0.135000 -0.060000 -0.04 ;
		RECT 0.060000 -0.135000 0.135000 -0.04 ;
		RECT -0.135000 0.060000 -0.060000 0.09 ;
		RECT 0.060000 0.060000 0.135000 0.09 ;
	LAYER M4 ;
		RECT -0.135000 -0.180000 0.135000 0.12 ;
END VIA34_4cut

VIA VIA34_FBD_XEN DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M3 ;
		RECT -0.037500 -0.037500 0.247500 0.085 ;
	LAYER VIA3 ;
		RECT 0.007500 0.007500 0.202500 0.055 ;
	LAYER M4 ;
		RECT -0.037500 -0.037500 0.247500 0.085 ;
END VIA34_FBD_XEN

VIA VIA34_FBD_XES DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M3 ;
		RECT -0.037500 -0.127500 0.247500 0.025 ;
	LAYER VIA3 ;
		RECT 0.007500 -0.082500 0.202500 -0.005 ;
	LAYER M4 ;
		RECT -0.037500 -0.127500 0.247500 0.025 ;
END VIA34_FBD_XES

VIA VIA34_FBD_XWN DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M3 ;
		RECT -0.247500 -0.037500 0.037500 0.085 ;
	LAYER VIA3 ;
		RECT -0.202500 0.007500 -0.007500 0.055 ;
	LAYER M4 ;
		RECT -0.247500 -0.037500 0.037500 0.085 ;
END VIA34_FBD_XWN

VIA VIA34_FBD_XWS DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M3 ;
		RECT -0.247500 -0.127500 0.037500 0.025 ;
	LAYER VIA3 ;
		RECT -0.202500 -0.082500 -0.007500 -0.005 ;
	LAYER M4 ;
		RECT -0.247500 -0.127500 0.037500 0.025 ;
END VIA34_FBD_XWS

VIA VIA34_FBD_YEN DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M3 ;
		RECT -0.037500 -0.037500 0.127500 0.165 ;
	LAYER VIA3 ;
		RECT 0.007500 0.007500 0.082500 0.135 ;
	LAYER M4 ;
		RECT -0.037500 -0.037500 0.127500 0.165 ;
END VIA34_FBD_YEN

VIA VIA34_FBD_YES DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M3 ;
		RECT -0.037500 -0.247500 0.127500 0.025 ;
	LAYER VIA3 ;
		RECT 0.007500 -0.202500 0.082500 -0.005 ;
	LAYER M4 ;
		RECT -0.037500 -0.247500 0.127500 0.025 ;
END VIA34_FBD_YES

VIA VIA34_FBD_YWN DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M3 ;
		RECT -0.127500 -0.037500 0.037500 0.165 ;
	LAYER VIA3 ;
		RECT -0.082500 0.007500 -0.007500 0.135 ;
	LAYER M4 ;
		RECT -0.127500 -0.037500 0.037500 0.165 ;
END VIA34_FBD_YWN

VIA VIA34_FBD_YWS DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M3 ;
		RECT -0.127500 -0.247500 0.037500 0.025 ;
	LAYER VIA3 ;
		RECT -0.082500 -0.202500 -0.007500 -0.005 ;
	LAYER M4 ;
		RECT -0.127500 -0.247500 0.037500 0.025 ;
END VIA34_FBD_YWS

VIA VIA34_FBS DEFAULT
	RESISTANCE 12.000000 ;
	LAYER M3 ;
		RECT -0.082500 -0.082500 0.082500 0.055 ;
	LAYER VIA3 ;
		RECT -0.037500 -0.037500 0.037500 0.025 ;
	LAYER M4 ;
		RECT -0.082500 -0.082500 0.082500 0.055 ;
END VIA34_FBS

VIA VIA34_FBS_EN DEFAULT
	RESISTANCE 12.000000 ;
	LAYER M3 ;
		RECT -0.037500 -0.037500 0.127500 0.085 ;
	LAYER VIA3 ;
		RECT 0.007500 0.007500 0.082500 0.055 ;
	LAYER M4 ;
		RECT -0.037500 -0.037500 0.127500 0.085 ;
END VIA34_FBS_EN

VIA VIA34_FBS_ES DEFAULT
	RESISTANCE 12.000000 ;
	LAYER M3 ;
		RECT -0.037500 -0.127500 0.127500 0.025 ;
	LAYER VIA3 ;
		RECT 0.007500 -0.082500 0.082500 -0.005 ;
	LAYER M4 ;
		RECT -0.037500 -0.127500 0.127500 0.025 ;
END VIA34_FBS_ES

VIA VIA34_FBS_WN DEFAULT
	RESISTANCE 12.000000 ;
	LAYER M3 ;
		RECT -0.127500 -0.037500 0.037500 0.085 ;
	LAYER VIA3 ;
		RECT -0.082500 0.007500 -0.007500 0.055 ;
	LAYER M4 ;
		RECT -0.127500 -0.037500 0.037500 0.085 ;
END VIA34_FBS_WN

VIA VIA34_FBS_WS DEFAULT
	RESISTANCE 12.000000 ;
	LAYER M3 ;
		RECT -0.127500 -0.127500 0.037500 0.025 ;
	LAYER VIA3 ;
		RECT -0.082500 -0.082500 -0.007500 -0.005 ;
	LAYER M4 ;
		RECT -0.127500 -0.127500 0.037500 0.025 ;
END VIA34_FBS_WS

VIA VIA34_PBD_E DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M3 ;
		RECT -0.052500 -0.037500 0.262500 0.025 ;
	LAYER VIA3 ;
		RECT 0.007500 -0.037500 0.202500 0.025 ;
	LAYER M4 ;
		RECT -0.037500 -0.082500 0.247500 0.055 ;
END VIA34_PBD_E

VIA VIA34_PBD_N DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M3 ;
		RECT -0.037500 -0.052500 0.037500 0.175 ;
	LAYER VIA3 ;
		RECT -0.037500 0.007500 0.037500 0.135 ;
	LAYER M4 ;
		RECT -0.082500 -0.037500 0.082500 0.165 ;
END VIA34_PBD_N

VIA VIA34_PBD_S DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M3 ;
		RECT -0.037500 -0.262500 0.037500 0.035 ;
	LAYER VIA3 ;
		RECT -0.037500 -0.202500 0.037500 -0.005 ;
	LAYER M4 ;
		RECT -0.082500 -0.247500 0.082500 0.025 ;
END VIA34_PBD_S

VIA VIA34_PBD_W DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M3 ;
		RECT -0.262500 -0.037500 0.052500 0.025 ;
	LAYER VIA3 ;
		RECT -0.202500 -0.037500 -0.007500 0.025 ;
	LAYER M4 ;
		RECT -0.247500 -0.082500 0.037500 0.055 ;
END VIA34_PBD_W

VIA VIA34_PBS_H DEFAULT
	RESISTANCE 12.000000 ;
	LAYER M3 ;
		RECT -0.082500 -0.037500 0.082500 0.025 ;
	LAYER VIA3 ;
		RECT -0.037500 -0.037500 0.037500 0.025 ;
	LAYER M4 ;
		RECT -0.082500 -0.082500 0.082500 0.055 ;
END VIA34_PBS_H

VIA VIA34_PBS_V DEFAULT
	RESISTANCE 12.000000 ;
	LAYER M3 ;
		RECT -0.037500 -0.082500 0.037500 0.055 ;
	LAYER VIA3 ;
		RECT -0.037500 -0.037500 0.037500 0.025 ;
	LAYER M4 ;
		RECT -0.082500 -0.082500 0.082500 0.055 ;
END VIA34_PBS_V

VIA VIA34_FBD20_XEN DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M3 ;
		RECT -0.037500 -0.037500 0.217500 0.065 ;
	LAYER VIA3 ;
		RECT -0.007500 -0.007500 0.187500 0.045 ;
	LAYER M4 ;
		RECT -0.037500 -0.037500 0.217500 0.065 ;
END VIA34_FBD20_XEN

VIA VIA34_FBD20_XES DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M3 ;
		RECT -0.037500 -0.097500 0.217500 0.025 ;
	LAYER VIA3 ;
		RECT -0.007500 -0.067500 0.187500 0.005 ;
	LAYER M4 ;
		RECT -0.037500 -0.097500 0.217500 0.025 ;
END VIA34_FBD20_XES

VIA VIA34_FBD20_XWN DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M3 ;
		RECT -0.217500 -0.037500 0.037500 0.065 ;
	LAYER VIA3 ;
		RECT -0.187500 -0.007500 0.007500 0.045 ;
	LAYER M4 ;
		RECT -0.217500 -0.037500 0.037500 0.065 ;
END VIA34_FBD20_XWN

VIA VIA34_FBD20_XWS DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M3 ;
		RECT -0.217500 -0.097500 0.037500 0.025 ;
	LAYER VIA3 ;
		RECT -0.187500 -0.067500 0.007500 0.005 ;
	LAYER M4 ;
		RECT -0.217500 -0.097500 0.037500 0.025 ;
END VIA34_FBD20_XWS

VIA VIA34_FBD20_YEN DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M3 ;
		RECT -0.037500 -0.037500 0.097500 0.145 ;
	LAYER VIA3 ;
		RECT -0.007500 -0.007500 0.067500 0.125 ;
	LAYER M4 ;
		RECT -0.037500 -0.037500 0.097500 0.145 ;
END VIA34_FBD20_YEN

VIA VIA34_FBD20_YES DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M3 ;
		RECT -0.037500 -0.217500 0.097500 0.025 ;
	LAYER VIA3 ;
		RECT -0.007500 -0.187500 0.067500 0.005 ;
	LAYER M4 ;
		RECT -0.037500 -0.217500 0.097500 0.025 ;
END VIA34_FBD20_YES

VIA VIA34_FBD20_YWN DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M3 ;
		RECT -0.097500 -0.037500 0.037500 0.145 ;
	LAYER VIA3 ;
		RECT -0.067500 -0.007500 0.007500 0.125 ;
	LAYER M4 ;
		RECT -0.097500 -0.037500 0.037500 0.145 ;
END VIA34_FBD20_YWN

VIA VIA34_FBD20_YWS DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M3 ;
		RECT -0.097500 -0.217500 0.037500 0.025 ;
	LAYER VIA3 ;
		RECT -0.067500 -0.187500 0.007500 0.005 ;
	LAYER M4 ;
		RECT -0.097500 -0.217500 0.037500 0.025 ;
END VIA34_FBD20_YWS

VIA VIA34_FBD30_XEN DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M3 ;
		RECT -0.037500 -0.037500 0.187500 0.085 ;
	LAYER VIA3 ;
		RECT -0.022500 0.007500 0.172500 0.055 ;
	LAYER M4 ;
		RECT -0.037500 -0.037500 0.187500 0.085 ;
END VIA34_FBD30_XEN

VIA VIA34_FBD30_XES DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M3 ;
		RECT -0.037500 -0.127500 0.187500 0.025 ;
	LAYER VIA3 ;
		RECT -0.022500 -0.082500 0.172500 -0.005 ;
	LAYER M4 ;
		RECT -0.037500 -0.127500 0.187500 0.025 ;
END VIA34_FBD30_XES

VIA VIA34_FBD30_XWN DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M3 ;
		RECT -0.187500 -0.037500 0.037500 0.085 ;
	LAYER VIA3 ;
		RECT -0.172500 0.007500 0.022500 0.055 ;
	LAYER M4 ;
		RECT -0.187500 -0.037500 0.037500 0.085 ;
END VIA34_FBD30_XWN

VIA VIA34_FBD30_XWS DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M3 ;
		RECT -0.187500 -0.127500 0.037500 0.025 ;
	LAYER VIA3 ;
		RECT -0.172500 -0.082500 0.022500 -0.005 ;
	LAYER M4 ;
		RECT -0.187500 -0.127500 0.037500 0.025 ;
END VIA34_FBD30_XWS

VIA VIA34_FBD30_YEN DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M3 ;
		RECT -0.037500 -0.037500 0.127500 0.125 ;
	LAYER VIA3 ;
		RECT 0.007500 -0.022500 0.082500 0.115 ;
	LAYER M4 ;
		RECT -0.037500 -0.037500 0.127500 0.125 ;
END VIA34_FBD30_YEN

VIA VIA34_FBD30_YES DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M3 ;
		RECT -0.037500 -0.187500 0.127500 0.025 ;
	LAYER VIA3 ;
		RECT 0.007500 -0.172500 0.082500 0.015 ;
	LAYER M4 ;
		RECT -0.037500 -0.187500 0.127500 0.025 ;
END VIA34_FBD30_YES

VIA VIA34_FBD30_YWN DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M3 ;
		RECT -0.127500 -0.037500 0.037500 0.125 ;
	LAYER VIA3 ;
		RECT -0.082500 -0.022500 -0.007500 0.115 ;
	LAYER M4 ;
		RECT -0.127500 -0.037500 0.037500 0.125 ;
END VIA34_FBD30_YWN

VIA VIA34_FBD30_YWS DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M3 ;
		RECT -0.127500 -0.187500 0.037500 0.025 ;
	LAYER VIA3 ;
		RECT -0.082500 -0.172500 -0.007500 0.015 ;
	LAYER M4 ;
		RECT -0.127500 -0.187500 0.037500 0.025 ;
END VIA34_FBD30_YWS

VIA VIA34_PBDB_E DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M3 ;
		RECT -0.007500 -0.067500 0.247500 0.045 ;
	LAYER VIA3 ;
		RECT 0.022500 -0.037500 0.217500 0.025 ;
	LAYER M4 ;
		RECT -0.037500 -0.037500 0.277500 0.025 ;
END VIA34_PBDB_E

VIA VIA34_PBDB_N DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M3 ;
		RECT -0.067500 -0.007500 0.067500 0.165 ;
	LAYER VIA3 ;
		RECT -0.037500 0.022500 0.037500 0.145 ;
	LAYER M4 ;
		RECT -0.037500 -0.037500 0.037500 0.185 ;
END VIA34_PBDB_N

VIA VIA34_PBDB_S DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M3 ;
		RECT -0.067500 -0.247500 0.067500 0.005 ;
	LAYER VIA3 ;
		RECT -0.037500 -0.217500 0.037500 -0.015 ;
	LAYER M4 ;
		RECT -0.037500 -0.277500 0.037500 0.025 ;
END VIA34_PBDB_S

VIA VIA34_PBDB_W DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M3 ;
		RECT -0.247500 -0.067500 0.007500 0.045 ;
	LAYER VIA3 ;
		RECT -0.217500 -0.037500 -0.022500 0.025 ;
	LAYER M4 ;
		RECT -0.277500 -0.037500 0.037500 0.025 ;
END VIA34_PBDB_W

VIA VIA34_PBDU_E DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M3 ;
		RECT -0.067500 -0.037500 0.247500 0.025 ;
	LAYER VIA3 ;
		RECT -0.007500 -0.037500 0.187500 0.025 ;
	LAYER M4 ;
		RECT -0.037500 -0.067500 0.217500 0.045 ;
END VIA34_PBDU_E

VIA VIA34_PBDU_N DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M3 ;
		RECT -0.037500 -0.067500 0.037500 0.165 ;
	LAYER VIA3 ;
		RECT -0.037500 -0.007500 0.037500 0.125 ;
	LAYER M4 ;
		RECT -0.067500 -0.037500 0.067500 0.145 ;
END VIA34_PBDU_N

VIA VIA34_PBDU_S DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M3 ;
		RECT -0.037500 -0.247500 0.037500 0.045 ;
	LAYER VIA3 ;
		RECT -0.037500 -0.187500 0.037500 0.005 ;
	LAYER M4 ;
		RECT -0.067500 -0.217500 0.067500 0.025 ;
END VIA34_PBDU_S

VIA VIA34_PBDU_W DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M3 ;
		RECT -0.247500 -0.037500 0.067500 0.025 ;
	LAYER VIA3 ;
		RECT -0.187500 -0.037500 0.007500 0.025 ;
	LAYER M4 ;
		RECT -0.217500 -0.067500 0.037500 0.045 ;
END VIA34_PBDU_W

VIA VIA34_PBDE_E DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M3 ;
		RECT -0.037500 -0.037500 0.277500 0.025 ;
	LAYER VIA3 ;
		RECT 0.022500 -0.037500 0.217500 0.025 ;
	LAYER M4 ;
		RECT -0.037500 -0.037500 0.277500 0.025 ;
END VIA34_PBDE_E

VIA VIA34_PBDE_N DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M3 ;
		RECT -0.037500 -0.037500 0.037500 0.185 ;
	LAYER VIA3 ;
		RECT -0.037500 0.022500 0.037500 0.145 ;
	LAYER M4 ;
		RECT -0.037500 -0.037500 0.037500 0.185 ;
END VIA34_PBDE_N

VIA VIA34_PBDE_S DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M3 ;
		RECT -0.037500 -0.277500 0.037500 0.025 ;
	LAYER VIA3 ;
		RECT -0.037500 -0.217500 0.037500 -0.015 ;
	LAYER M4 ;
		RECT -0.037500 -0.277500 0.037500 0.025 ;
END VIA34_PBDE_S

VIA VIA34_PBDE_W DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M3 ;
		RECT -0.277500 -0.037500 0.037500 0.025 ;
	LAYER VIA3 ;
		RECT -0.217500 -0.037500 -0.022500 0.025 ;
	LAYER M4 ;
		RECT -0.277500 -0.037500 0.037500 0.025 ;
END VIA34_PBDE_W

VIA VIA34_FBS25 DEFAULT
	RESISTANCE 12.000000 ;
	LAYER M3 ;
		RECT -0.075000 -0.075000 0.075000 0.05 ;
	LAYER VIA3 ;
		RECT -0.037500 -0.037500 0.037500 0.025 ;
	LAYER M4 ;
		RECT -0.075000 -0.075000 0.075000 0.05 ;
END VIA34_FBS25

VIA VIA34_FBS25_EN DEFAULT
	RESISTANCE 12.000000 ;
	LAYER M3 ;
		RECT -0.037500 -0.037500 0.112500 0.075 ;
	LAYER VIA3 ;
		RECT 0.000000 0.000000 0.075000 0.05 ;
	LAYER M4 ;
		RECT -0.037500 -0.037500 0.112500 0.075 ;
END VIA34_FBS25_EN

VIA VIA34_FBS25_ES DEFAULT
	RESISTANCE 12.000000 ;
	LAYER M3 ;
		RECT -0.037500 -0.112500 0.112500 0.025 ;
	LAYER VIA3 ;
		RECT 0.000000 -0.075000 0.075000 0 ;
	LAYER M4 ;
		RECT -0.037500 -0.112500 0.112500 0.025 ;
END VIA34_FBS25_ES

VIA VIA34_FBS25_WN DEFAULT
	RESISTANCE 12.000000 ;
	LAYER M3 ;
		RECT -0.112500 -0.037500 0.037500 0.075 ;
	LAYER VIA3 ;
		RECT -0.075000 0.000000 0.000000 0.05 ;
	LAYER M4 ;
		RECT -0.112500 -0.037500 0.037500 0.075 ;
END VIA34_FBS25_WN

VIA VIA34_FBS25_WS DEFAULT
	RESISTANCE 12.000000 ;
	LAYER M3 ;
		RECT -0.112500 -0.112500 0.037500 0.025 ;
	LAYER VIA3 ;
		RECT -0.075000 -0.075000 0.000000 0 ;
	LAYER M4 ;
		RECT -0.112500 -0.112500 0.037500 0.025 ;
END VIA34_FBS25_WS

VIA VIA34_PBSU_H DEFAULT
	RESISTANCE 12.000000 ;
	LAYER M3 ;
		RECT -0.082500 -0.037500 0.082500 0.025 ;
	LAYER VIA3 ;
		RECT -0.037500 -0.037500 0.037500 0.025 ;
	LAYER M4 ;
		RECT -0.052500 -0.075000 0.052500 0.05 ;
END VIA34_PBSU_H

VIA VIA34_PBSU_V DEFAULT
	RESISTANCE 12.000000 ;
	LAYER M3 ;
		RECT -0.037500 -0.082500 0.037500 0.055 ;
	LAYER VIA3 ;
		RECT -0.037500 -0.037500 0.037500 0.025 ;
	LAYER M4 ;
		RECT -0.075000 -0.052500 0.075000 0.035 ;
END VIA34_PBSU_V

VIA VIA34_PBSB_H DEFAULT
	RESISTANCE 12.000000 ;
	LAYER M3 ;
		RECT -0.075000 -0.052500 0.075000 0.035 ;
	LAYER VIA3 ;
		RECT -0.037500 -0.037500 0.037500 0.025 ;
	LAYER M4 ;
		RECT -0.037500 -0.082500 0.037500 0.055 ;
END VIA34_PBSB_H

VIA VIA34_PBSB_V DEFAULT
	RESISTANCE 12.000000 ;
	LAYER M3 ;
		RECT -0.052500 -0.075000 0.052500 0.05 ;
	LAYER VIA3 ;
		RECT -0.037500 -0.037500 0.037500 0.025 ;
	LAYER M4 ;
		RECT -0.082500 -0.037500 0.082500 0.025 ;
END VIA34_PBSB_V


VIA VIA45_1cut DEFAULT
	RESISTANCE 12.000000 ;
	LAYER M4 ;
		RECT -0.037500 -0.082500 0.037500 0.055 ;
	LAYER VIA4 ;
		RECT -0.037500 -0.037500 0.037500 0.025 ;
	LAYER M5 ;
		RECT -0.082500 -0.037500 0.082500 0.025 ;
END VIA45_1cut

VIA VIA45_1cut_FAT_C DEFAULT
	RESISTANCE 12.000000 ;
	LAYER M4 ;
		RECT -0.037500 -0.112500 0.037500 0.075 ;
	LAYER VIA4 ;
		RECT -0.037500 -0.037500 0.037500 0.025 ;
	LAYER M5 ;
		RECT -0.112500 -0.037500 0.112500 0.025 ;
END VIA45_1cut_FAT_C

VIA VIA45_1cut_EN1415 DEFAULT
	RESISTANCE 12.000000 ;
	LAYER M4 ;
		RECT -0.052500 -0.075000 0.052500 0.05 ;
	LAYER VIA4 ;
		RECT -0.037500 -0.037500 0.037500 0.025 ;
	LAYER M5 ;
		RECT -0.075000 -0.052500 0.075000 0.035 ;
END VIA45_1cut_EN1415

VIA VIA45_1stack_C DEFAULT
	RESISTANCE 12.000000 ;
	LAYER M4 ;
		RECT -0.037500 -0.255000 0.037500 0.17 ;
	LAYER VIA4 ;
		RECT -0.037500 -0.037500 0.037500 0.025 ;
	LAYER M5 ;
		RECT -0.082500 -0.037500 0.082500 0.025 ;
END VIA45_1stack_C

VIA VIA45_1stack_N DEFAULT
	RESISTANCE 12.000000 ;
	LAYER M4 ;
		RECT -0.037500 -0.082500 0.037500 0.285 ;
	LAYER VIA4 ;
		RECT -0.037500 -0.037500 0.037500 0.025 ;
	LAYER M5 ;
		RECT -0.082500 -0.037500 0.082500 0.025 ;
END VIA45_1stack_N

VIA VIA45_1stack_S DEFAULT
	RESISTANCE 12.000000 ;
	LAYER M4 ;
		RECT -0.037500 -0.427500 0.037500 0.055 ;
	LAYER VIA4 ;
		RECT -0.037500 -0.037500 0.037500 0.025 ;
	LAYER M5 ;
		RECT -0.082500 -0.037500 0.082500 0.025 ;
END VIA45_1stack_S

VIA VIA45_2cut_P1_N DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M4 ;
		RECT -0.037500 -0.082500 0.037500 0.155 ;
	LAYER VIA4 ;
		RECT -0.037500 -0.022500 0.037500 0.115 ;
	LAYER M5 ;
		RECT -0.082500 -0.037500 0.082500 0.125 ;
END VIA45_2cut_P1_N

VIA VIA45_2cut_P1_S DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M4 ;
		RECT -0.037500 -0.232500 0.037500 0.055 ;
	LAYER VIA4 ;
		RECT -0.037500 -0.172500 0.037500 0.015 ;
	LAYER M5 ;
		RECT -0.082500 -0.187500 0.082500 0.025 ;
END VIA45_2cut_P1_S

VIA VIA45_2cut_P2_BLC DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M4 ;
		RECT -0.112500 -0.082500 0.112500 0.055 ;
	LAYER VIA4 ;
		RECT -0.097500 -0.037500 0.097500 0.025 ;
	LAYER M5 ;
		RECT -0.330000 -0.037500 0.330000 0.025 ;
END VIA45_2cut_P2_BLC

VIA VIA45_2cut_P2_BLE DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M4 ;
		RECT -0.037500 -0.082500 0.187500 0.055 ;
	LAYER VIA4 ;
		RECT -0.022500 -0.037500 0.172500 0.025 ;
	LAYER M5 ;
		RECT -0.255000 -0.037500 0.405000 0.025 ;
END VIA45_2cut_P2_BLE

VIA VIA45_2cut_P2_BLW DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M4 ;
		RECT -0.187500 -0.082500 0.037500 0.055 ;
	LAYER VIA4 ;
		RECT -0.172500 -0.037500 0.022500 0.025 ;
	LAYER M5 ;
		RECT -0.405000 -0.037500 0.255000 0.025 ;
END VIA45_2cut_P2_BLW

VIA VIA45_2cut_P2_SLE DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M4 ;
		RECT -0.037500 -0.082500 0.187500 0.055 ;
	LAYER VIA4 ;
		RECT -0.022500 -0.037500 0.172500 0.025 ;
	LAYER M5 ;
		RECT -0.097500 -0.037500 0.562500 0.025 ;
END VIA45_2cut_P2_SLE

VIA VIA45_2cut_P2_SLW DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M4 ;
		RECT -0.187500 -0.082500 0.037500 0.055 ;
	LAYER VIA4 ;
		RECT -0.172500 -0.037500 0.022500 0.025 ;
	LAYER M5 ;
		RECT -0.562500 -0.037500 0.097500 0.025 ;
END VIA45_2cut_P2_SLW

VIA VIA45_2cut_P3_E DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M4 ;
		RECT -0.037500 -0.082500 0.187500 0.055 ;
	LAYER VIA4 ;
		RECT -0.022500 -0.037500 0.172500 0.025 ;
	LAYER M5 ;
		RECT -0.082500 -0.037500 0.232500 0.025 ;
END VIA45_2cut_P3_E

VIA VIA45_2cut_P3_W DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M4 ;
		RECT -0.187500 -0.082500 0.037500 0.055 ;
	LAYER VIA4 ;
		RECT -0.172500 -0.037500 0.022500 0.025 ;
	LAYER M5 ;
		RECT -0.232500 -0.037500 0.082500 0.025 ;
END VIA45_2cut_P3_W

VIA VIA45_4cut DEFAULT
	RESISTANCE 3.000000 ;
	LAYER M4 ;
		RECT -0.135000 -0.180000 0.135000 0.12 ;
	LAYER VIA4 ;
		RECT -0.135000 -0.135000 -0.060000 -0.04 ;
		RECT 0.060000 -0.135000 0.135000 -0.04 ;
		RECT -0.135000 0.060000 -0.060000 0.09 ;
		RECT 0.060000 0.060000 0.135000 0.09 ;
	LAYER M5 ;
		RECT -0.180000 -0.135000 0.180000 0.09 ;
END VIA45_4cut

VIA VIA45_FBD_XEN DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M4 ;
		RECT -0.037500 -0.037500 0.247500 0.085 ;
	LAYER VIA4 ;
		RECT 0.007500 0.007500 0.202500 0.055 ;
	LAYER M5 ;
		RECT -0.037500 -0.037500 0.247500 0.085 ;
END VIA45_FBD_XEN

VIA VIA45_FBD_XES DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M4 ;
		RECT -0.037500 -0.127500 0.247500 0.025 ;
	LAYER VIA4 ;
		RECT 0.007500 -0.082500 0.202500 -0.005 ;
	LAYER M5 ;
		RECT -0.037500 -0.127500 0.247500 0.025 ;
END VIA45_FBD_XES

VIA VIA45_FBD_XWN DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M4 ;
		RECT -0.247500 -0.037500 0.037500 0.085 ;
	LAYER VIA4 ;
		RECT -0.202500 0.007500 -0.007500 0.055 ;
	LAYER M5 ;
		RECT -0.247500 -0.037500 0.037500 0.085 ;
END VIA45_FBD_XWN

VIA VIA45_FBD_XWS DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M4 ;
		RECT -0.247500 -0.127500 0.037500 0.025 ;
	LAYER VIA4 ;
		RECT -0.202500 -0.082500 -0.007500 -0.005 ;
	LAYER M5 ;
		RECT -0.247500 -0.127500 0.037500 0.025 ;
END VIA45_FBD_XWS

VIA VIA45_FBD_YEN DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M4 ;
		RECT -0.037500 -0.037500 0.127500 0.165 ;
	LAYER VIA4 ;
		RECT 0.007500 0.007500 0.082500 0.135 ;
	LAYER M5 ;
		RECT -0.037500 -0.037500 0.127500 0.165 ;
END VIA45_FBD_YEN

VIA VIA45_FBD_YES DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M4 ;
		RECT -0.037500 -0.247500 0.127500 0.025 ;
	LAYER VIA4 ;
		RECT 0.007500 -0.202500 0.082500 -0.005 ;
	LAYER M5 ;
		RECT -0.037500 -0.247500 0.127500 0.025 ;
END VIA45_FBD_YES

VIA VIA45_FBD_YWN DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M4 ;
		RECT -0.127500 -0.037500 0.037500 0.165 ;
	LAYER VIA4 ;
		RECT -0.082500 0.007500 -0.007500 0.135 ;
	LAYER M5 ;
		RECT -0.127500 -0.037500 0.037500 0.165 ;
END VIA45_FBD_YWN

VIA VIA45_FBD_YWS DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M4 ;
		RECT -0.127500 -0.247500 0.037500 0.025 ;
	LAYER VIA4 ;
		RECT -0.082500 -0.202500 -0.007500 -0.005 ;
	LAYER M5 ;
		RECT -0.127500 -0.247500 0.037500 0.025 ;
END VIA45_FBD_YWS

VIA VIA45_FBS DEFAULT
	RESISTANCE 12.000000 ;
	LAYER M4 ;
		RECT -0.082500 -0.082500 0.082500 0.055 ;
	LAYER VIA4 ;
		RECT -0.037500 -0.037500 0.037500 0.025 ;
	LAYER M5 ;
		RECT -0.082500 -0.082500 0.082500 0.055 ;
END VIA45_FBS

VIA VIA45_FBS_EN DEFAULT
	RESISTANCE 12.000000 ;
	LAYER M4 ;
		RECT -0.037500 -0.037500 0.127500 0.085 ;
	LAYER VIA4 ;
		RECT 0.007500 0.007500 0.082500 0.055 ;
	LAYER M5 ;
		RECT -0.037500 -0.037500 0.127500 0.085 ;
END VIA45_FBS_EN

VIA VIA45_FBS_ES DEFAULT
	RESISTANCE 12.000000 ;
	LAYER M4 ;
		RECT -0.037500 -0.127500 0.127500 0.025 ;
	LAYER VIA4 ;
		RECT 0.007500 -0.082500 0.082500 -0.005 ;
	LAYER M5 ;
		RECT -0.037500 -0.127500 0.127500 0.025 ;
END VIA45_FBS_ES

VIA VIA45_FBS_WN DEFAULT
	RESISTANCE 12.000000 ;
	LAYER M4 ;
		RECT -0.127500 -0.037500 0.037500 0.085 ;
	LAYER VIA4 ;
		RECT -0.082500 0.007500 -0.007500 0.055 ;
	LAYER M5 ;
		RECT -0.127500 -0.037500 0.037500 0.085 ;
END VIA45_FBS_WN

VIA VIA45_FBS_WS DEFAULT
	RESISTANCE 12.000000 ;
	LAYER M4 ;
		RECT -0.127500 -0.127500 0.037500 0.025 ;
	LAYER VIA4 ;
		RECT -0.082500 -0.082500 -0.007500 -0.005 ;
	LAYER M5 ;
		RECT -0.127500 -0.127500 0.037500 0.025 ;
END VIA45_FBS_WS

VIA VIA45_PBD_E DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M4 ;
		RECT -0.052500 -0.037500 0.262500 0.025 ;
	LAYER VIA4 ;
		RECT 0.007500 -0.037500 0.202500 0.025 ;
	LAYER M5 ;
		RECT -0.037500 -0.082500 0.247500 0.055 ;
END VIA45_PBD_E

VIA VIA45_PBD_N DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M4 ;
		RECT -0.037500 -0.052500 0.037500 0.175 ;
	LAYER VIA4 ;
		RECT -0.037500 0.007500 0.037500 0.135 ;
	LAYER M5 ;
		RECT -0.082500 -0.037500 0.082500 0.165 ;
END VIA45_PBD_N

VIA VIA45_PBD_S DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M4 ;
		RECT -0.037500 -0.262500 0.037500 0.035 ;
	LAYER VIA4 ;
		RECT -0.037500 -0.202500 0.037500 -0.005 ;
	LAYER M5 ;
		RECT -0.082500 -0.247500 0.082500 0.025 ;
END VIA45_PBD_S

VIA VIA45_PBD_W DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M4 ;
		RECT -0.262500 -0.037500 0.052500 0.025 ;
	LAYER VIA4 ;
		RECT -0.202500 -0.037500 -0.007500 0.025 ;
	LAYER M5 ;
		RECT -0.247500 -0.082500 0.037500 0.055 ;
END VIA45_PBD_W

VIA VIA45_PBS_H DEFAULT
	RESISTANCE 12.000000 ;
	LAYER M4 ;
		RECT -0.082500 -0.037500 0.082500 0.025 ;
	LAYER VIA4 ;
		RECT -0.037500 -0.037500 0.037500 0.025 ;
	LAYER M5 ;
		RECT -0.082500 -0.082500 0.082500 0.055 ;
END VIA45_PBS_H

VIA VIA45_PBS_V DEFAULT
	RESISTANCE 12.000000 ;
	LAYER M4 ;
		RECT -0.037500 -0.082500 0.037500 0.055 ;
	LAYER VIA4 ;
		RECT -0.037500 -0.037500 0.037500 0.025 ;
	LAYER M5 ;
		RECT -0.082500 -0.082500 0.082500 0.055 ;
END VIA45_PBS_V

VIA VIA45_FBD20_XEN DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M4 ;
		RECT -0.037500 -0.037500 0.217500 0.065 ;
	LAYER VIA4 ;
		RECT -0.007500 -0.007500 0.187500 0.045 ;
	LAYER M5 ;
		RECT -0.037500 -0.037500 0.217500 0.065 ;
END VIA45_FBD20_XEN

VIA VIA45_FBD20_XES DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M4 ;
		RECT -0.037500 -0.097500 0.217500 0.025 ;
	LAYER VIA4 ;
		RECT -0.007500 -0.067500 0.187500 0.005 ;
	LAYER M5 ;
		RECT -0.037500 -0.097500 0.217500 0.025 ;
END VIA45_FBD20_XES

VIA VIA45_FBD20_XWN DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M4 ;
		RECT -0.217500 -0.037500 0.037500 0.065 ;
	LAYER VIA4 ;
		RECT -0.187500 -0.007500 0.007500 0.045 ;
	LAYER M5 ;
		RECT -0.217500 -0.037500 0.037500 0.065 ;
END VIA45_FBD20_XWN

VIA VIA45_FBD20_XWS DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M4 ;
		RECT -0.217500 -0.097500 0.037500 0.025 ;
	LAYER VIA4 ;
		RECT -0.187500 -0.067500 0.007500 0.005 ;
	LAYER M5 ;
		RECT -0.217500 -0.097500 0.037500 0.025 ;
END VIA45_FBD20_XWS

VIA VIA45_FBD20_YEN DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M4 ;
		RECT -0.037500 -0.037500 0.097500 0.145 ;
	LAYER VIA4 ;
		RECT -0.007500 -0.007500 0.067500 0.125 ;
	LAYER M5 ;
		RECT -0.037500 -0.037500 0.097500 0.145 ;
END VIA45_FBD20_YEN

VIA VIA45_FBD20_YES DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M4 ;
		RECT -0.037500 -0.217500 0.097500 0.025 ;
	LAYER VIA4 ;
		RECT -0.007500 -0.187500 0.067500 0.005 ;
	LAYER M5 ;
		RECT -0.037500 -0.217500 0.097500 0.025 ;
END VIA45_FBD20_YES

VIA VIA45_FBD20_YWN DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M4 ;
		RECT -0.097500 -0.037500 0.037500 0.145 ;
	LAYER VIA4 ;
		RECT -0.067500 -0.007500 0.007500 0.125 ;
	LAYER M5 ;
		RECT -0.097500 -0.037500 0.037500 0.145 ;
END VIA45_FBD20_YWN

VIA VIA45_FBD20_YWS DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M4 ;
		RECT -0.097500 -0.217500 0.037500 0.025 ;
	LAYER VIA4 ;
		RECT -0.067500 -0.187500 0.007500 0.005 ;
	LAYER M5 ;
		RECT -0.097500 -0.217500 0.037500 0.025 ;
END VIA45_FBD20_YWS

VIA VIA45_FBD30_XEN DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M4 ;
		RECT -0.037500 -0.037500 0.187500 0.085 ;
	LAYER VIA4 ;
		RECT -0.022500 0.007500 0.172500 0.055 ;
	LAYER M5 ;
		RECT -0.037500 -0.037500 0.187500 0.085 ;
END VIA45_FBD30_XEN

VIA VIA45_FBD30_XES DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M4 ;
		RECT -0.037500 -0.127500 0.187500 0.025 ;
	LAYER VIA4 ;
		RECT -0.022500 -0.082500 0.172500 -0.005 ;
	LAYER M5 ;
		RECT -0.037500 -0.127500 0.187500 0.025 ;
END VIA45_FBD30_XES

VIA VIA45_FBD30_XWN DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M4 ;
		RECT -0.187500 -0.037500 0.037500 0.085 ;
	LAYER VIA4 ;
		RECT -0.172500 0.007500 0.022500 0.055 ;
	LAYER M5 ;
		RECT -0.187500 -0.037500 0.037500 0.085 ;
END VIA45_FBD30_XWN

VIA VIA45_FBD30_XWS DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M4 ;
		RECT -0.187500 -0.127500 0.037500 0.025 ;
	LAYER VIA4 ;
		RECT -0.172500 -0.082500 0.022500 -0.005 ;
	LAYER M5 ;
		RECT -0.187500 -0.127500 0.037500 0.025 ;
END VIA45_FBD30_XWS

VIA VIA45_FBD30_YEN DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M4 ;
		RECT -0.037500 -0.037500 0.127500 0.125 ;
	LAYER VIA4 ;
		RECT 0.007500 -0.022500 0.082500 0.115 ;
	LAYER M5 ;
		RECT -0.037500 -0.037500 0.127500 0.125 ;
END VIA45_FBD30_YEN

VIA VIA45_FBD30_YES DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M4 ;
		RECT -0.037500 -0.187500 0.127500 0.025 ;
	LAYER VIA4 ;
		RECT 0.007500 -0.172500 0.082500 0.015 ;
	LAYER M5 ;
		RECT -0.037500 -0.187500 0.127500 0.025 ;
END VIA45_FBD30_YES

VIA VIA45_FBD30_YWN DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M4 ;
		RECT -0.127500 -0.037500 0.037500 0.125 ;
	LAYER VIA4 ;
		RECT -0.082500 -0.022500 -0.007500 0.115 ;
	LAYER M5 ;
		RECT -0.127500 -0.037500 0.037500 0.125 ;
END VIA45_FBD30_YWN

VIA VIA45_FBD30_YWS DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M4 ;
		RECT -0.127500 -0.187500 0.037500 0.025 ;
	LAYER VIA4 ;
		RECT -0.082500 -0.172500 -0.007500 0.015 ;
	LAYER M5 ;
		RECT -0.127500 -0.187500 0.037500 0.025 ;
END VIA45_FBD30_YWS

VIA VIA45_PBDB_E DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M4 ;
		RECT -0.007500 -0.067500 0.247500 0.045 ;
	LAYER VIA4 ;
		RECT 0.022500 -0.037500 0.217500 0.025 ;
	LAYER M5 ;
		RECT -0.037500 -0.037500 0.277500 0.025 ;
END VIA45_PBDB_E

VIA VIA45_PBDB_N DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M4 ;
		RECT -0.067500 -0.007500 0.067500 0.165 ;
	LAYER VIA4 ;
		RECT -0.037500 0.022500 0.037500 0.145 ;
	LAYER M5 ;
		RECT -0.037500 -0.037500 0.037500 0.185 ;
END VIA45_PBDB_N

VIA VIA45_PBDB_S DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M4 ;
		RECT -0.067500 -0.247500 0.067500 0.005 ;
	LAYER VIA4 ;
		RECT -0.037500 -0.217500 0.037500 -0.015 ;
	LAYER M5 ;
		RECT -0.037500 -0.277500 0.037500 0.025 ;
END VIA45_PBDB_S

VIA VIA45_PBDB_W DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M4 ;
		RECT -0.247500 -0.067500 0.007500 0.045 ;
	LAYER VIA4 ;
		RECT -0.217500 -0.037500 -0.022500 0.025 ;
	LAYER M5 ;
		RECT -0.277500 -0.037500 0.037500 0.025 ;
END VIA45_PBDB_W

VIA VIA45_PBDU_E DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M4 ;
		RECT -0.067500 -0.037500 0.247500 0.025 ;
	LAYER VIA4 ;
		RECT -0.007500 -0.037500 0.187500 0.025 ;
	LAYER M5 ;
		RECT -0.037500 -0.067500 0.217500 0.045 ;
END VIA45_PBDU_E

VIA VIA45_PBDU_N DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M4 ;
		RECT -0.037500 -0.067500 0.037500 0.165 ;
	LAYER VIA4 ;
		RECT -0.037500 -0.007500 0.037500 0.125 ;
	LAYER M5 ;
		RECT -0.067500 -0.037500 0.067500 0.145 ;
END VIA45_PBDU_N

VIA VIA45_PBDU_S DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M4 ;
		RECT -0.037500 -0.247500 0.037500 0.045 ;
	LAYER VIA4 ;
		RECT -0.037500 -0.187500 0.037500 0.005 ;
	LAYER M5 ;
		RECT -0.067500 -0.217500 0.067500 0.025 ;
END VIA45_PBDU_S

VIA VIA45_PBDU_W DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M4 ;
		RECT -0.247500 -0.037500 0.067500 0.025 ;
	LAYER VIA4 ;
		RECT -0.187500 -0.037500 0.007500 0.025 ;
	LAYER M5 ;
		RECT -0.217500 -0.067500 0.037500 0.045 ;
END VIA45_PBDU_W

VIA VIA45_PBDE_E DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M4 ;
		RECT -0.037500 -0.037500 0.277500 0.025 ;
	LAYER VIA4 ;
		RECT 0.022500 -0.037500 0.217500 0.025 ;
	LAYER M5 ;
		RECT -0.037500 -0.037500 0.277500 0.025 ;
END VIA45_PBDE_E

VIA VIA45_PBDE_N DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M4 ;
		RECT -0.037500 -0.037500 0.037500 0.185 ;
	LAYER VIA4 ;
		RECT -0.037500 0.022500 0.037500 0.145 ;
	LAYER M5 ;
		RECT -0.037500 -0.037500 0.037500 0.185 ;
END VIA45_PBDE_N

VIA VIA45_PBDE_S DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M4 ;
		RECT -0.037500 -0.277500 0.037500 0.025 ;
	LAYER VIA4 ;
		RECT -0.037500 -0.217500 0.037500 -0.015 ;
	LAYER M5 ;
		RECT -0.037500 -0.277500 0.037500 0.025 ;
END VIA45_PBDE_S

VIA VIA45_PBDE_W DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M4 ;
		RECT -0.277500 -0.037500 0.037500 0.025 ;
	LAYER VIA4 ;
		RECT -0.217500 -0.037500 -0.022500 0.025 ;
	LAYER M5 ;
		RECT -0.277500 -0.037500 0.037500 0.025 ;
END VIA45_PBDE_W

VIA VIA45_FBS25 DEFAULT
	RESISTANCE 12.000000 ;
	LAYER M4 ;
		RECT -0.075000 -0.075000 0.075000 0.05 ;
	LAYER VIA4 ;
		RECT -0.037500 -0.037500 0.037500 0.025 ;
	LAYER M5 ;
		RECT -0.075000 -0.075000 0.075000 0.05 ;
END VIA45_FBS25

VIA VIA45_FBS25_EN DEFAULT
	RESISTANCE 12.000000 ;
	LAYER M4 ;
		RECT -0.037500 -0.037500 0.112500 0.075 ;
	LAYER VIA4 ;
		RECT 0.000000 0.000000 0.075000 0.05 ;
	LAYER M5 ;
		RECT -0.037500 -0.037500 0.112500 0.075 ;
END VIA45_FBS25_EN

VIA VIA45_FBS25_ES DEFAULT
	RESISTANCE 12.000000 ;
	LAYER M4 ;
		RECT -0.037500 -0.112500 0.112500 0.025 ;
	LAYER VIA4 ;
		RECT 0.000000 -0.075000 0.075000 0 ;
	LAYER M5 ;
		RECT -0.037500 -0.112500 0.112500 0.025 ;
END VIA45_FBS25_ES

VIA VIA45_FBS25_WN DEFAULT
	RESISTANCE 12.000000 ;
	LAYER M4 ;
		RECT -0.112500 -0.037500 0.037500 0.075 ;
	LAYER VIA4 ;
		RECT -0.075000 0.000000 0.000000 0.05 ;
	LAYER M5 ;
		RECT -0.112500 -0.037500 0.037500 0.075 ;
END VIA45_FBS25_WN

VIA VIA45_FBS25_WS DEFAULT
	RESISTANCE 12.000000 ;
	LAYER M4 ;
		RECT -0.112500 -0.112500 0.037500 0.025 ;
	LAYER VIA4 ;
		RECT -0.075000 -0.075000 0.000000 0 ;
	LAYER M5 ;
		RECT -0.112500 -0.112500 0.037500 0.025 ;
END VIA45_FBS25_WS

VIA VIA45_PBSU_H DEFAULT
	RESISTANCE 12.000000 ;
	LAYER M4 ;
		RECT -0.082500 -0.037500 0.082500 0.025 ;
	LAYER VIA4 ;
		RECT -0.037500 -0.037500 0.037500 0.025 ;
	LAYER M5 ;
		RECT -0.052500 -0.075000 0.052500 0.05 ;
END VIA45_PBSU_H

VIA VIA45_PBSU_V DEFAULT
	RESISTANCE 12.000000 ;
	LAYER M4 ;
		RECT -0.037500 -0.082500 0.037500 0.055 ;
	LAYER VIA4 ;
		RECT -0.037500 -0.037500 0.037500 0.025 ;
	LAYER M5 ;
		RECT -0.075000 -0.052500 0.075000 0.035 ;
END VIA45_PBSU_V

VIA VIA45_PBSB_H DEFAULT
	RESISTANCE 12.000000 ;
	LAYER M4 ;
		RECT -0.075000 -0.052500 0.075000 0.035 ;
	LAYER VIA4 ;
		RECT -0.037500 -0.037500 0.037500 0.025 ;
	LAYER M5 ;
		RECT -0.037500 -0.082500 0.037500 0.055 ;
END VIA45_PBSB_H

VIA VIA45_PBSB_V DEFAULT
	RESISTANCE 12.000000 ;
	LAYER M4 ;
		RECT -0.052500 -0.075000 0.052500 0.05 ;
	LAYER VIA4 ;
		RECT -0.037500 -0.037500 0.037500 0.025 ;
	LAYER M5 ;
		RECT -0.082500 -0.037500 0.082500 0.025 ;
END VIA45_PBSB_V


VIA VIA56_1cut DEFAULT
	RESISTANCE 12.000000 ;
	LAYER M5 ;
		RECT -0.082500 -0.037500 0.082500 0.025 ;
	LAYER VIA5 ;
		RECT -0.037500 -0.037500 0.037500 0.025 ;
	LAYER M6 ;
		RECT -0.037500 -0.082500 0.037500 0.055 ;
END VIA56_1cut

VIA VIA56_1cut_FAT_C DEFAULT
	RESISTANCE 12.000000 ;
	LAYER M5 ;
		RECT -0.112500 -0.037500 0.112500 0.025 ;
	LAYER VIA5 ;
		RECT -0.037500 -0.037500 0.037500 0.025 ;
	LAYER M6 ;
		RECT -0.037500 -0.112500 0.037500 0.075 ;
END VIA56_1cut_FAT_C

VIA VIA56_1cut_EN1415 DEFAULT
	RESISTANCE 12.000000 ;
	LAYER M5 ;
		RECT -0.075000 -0.052500 0.075000 0.035 ;
	LAYER VIA5 ;
		RECT -0.037500 -0.037500 0.037500 0.025 ;
	LAYER M6 ;
		RECT -0.052500 -0.075000 0.052500 0.05 ;
END VIA56_1cut_EN1415

VIA VIA56_1stack_C DEFAULT
	RESISTANCE 12.000000 ;
	LAYER M5 ;
		RECT -0.255000 -0.037500 0.255000 0.025 ;
	LAYER VIA5 ;
		RECT -0.037500 -0.037500 0.037500 0.025 ;
	LAYER M6 ;
		RECT -0.037500 -0.082500 0.037500 0.055 ;
END VIA56_1stack_C

VIA VIA56_1stack_E DEFAULT
	RESISTANCE 12.000000 ;
	LAYER M5 ;
		RECT -0.082500 -0.037500 0.427500 0.025 ;
	LAYER VIA5 ;
		RECT -0.037500 -0.037500 0.037500 0.025 ;
	LAYER M6 ;
		RECT -0.037500 -0.082500 0.037500 0.055 ;
END VIA56_1stack_E

VIA VIA56_1stack_W DEFAULT
	RESISTANCE 12.000000 ;
	LAYER M5 ;
		RECT -0.427500 -0.037500 0.082500 0.025 ;
	LAYER VIA5 ;
		RECT -0.037500 -0.037500 0.037500 0.025 ;
	LAYER M6 ;
		RECT -0.037500 -0.082500 0.037500 0.055 ;
END VIA56_1stack_W

VIA VIA56_2cut_P1_E DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M5 ;
		RECT -0.082500 -0.037500 0.232500 0.025 ;
	LAYER VIA5 ;
		RECT -0.022500 -0.037500 0.172500 0.025 ;
	LAYER M6 ;
		RECT -0.037500 -0.082500 0.187500 0.055 ;
END VIA56_2cut_P1_E

VIA VIA56_2cut_P1_W DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M5 ;
		RECT -0.232500 -0.037500 0.082500 0.025 ;
	LAYER VIA5 ;
		RECT -0.172500 -0.037500 0.022500 0.025 ;
	LAYER M6 ;
		RECT -0.187500 -0.082500 0.037500 0.055 ;
END VIA56_2cut_P1_W

VIA VIA56_2cut_P2_BLC DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M5 ;
		RECT -0.082500 -0.112500 0.082500 0.075 ;
	LAYER VIA5 ;
		RECT -0.037500 -0.097500 0.037500 0.065 ;
	LAYER M6 ;
		RECT -0.037500 -0.330000 0.037500 0.22 ;
END VIA56_2cut_P2_BLC

VIA VIA56_2cut_P2_BLN DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M5 ;
		RECT -0.082500 -0.037500 0.082500 0.125 ;
	LAYER VIA5 ;
		RECT -0.037500 -0.022500 0.037500 0.115 ;
	LAYER M6 ;
		RECT -0.037500 -0.255000 0.037500 0.27 ;
END VIA56_2cut_P2_BLN

VIA VIA56_2cut_P2_BLS DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M5 ;
		RECT -0.082500 -0.187500 0.082500 0.025 ;
	LAYER VIA5 ;
		RECT -0.037500 -0.172500 0.037500 0.015 ;
	LAYER M6 ;
		RECT -0.037500 -0.405000 0.037500 0.17 ;
END VIA56_2cut_P2_BLS

VIA VIA56_2cut_P2_SLN DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M5 ;
		RECT -0.082500 -0.037500 0.082500 0.125 ;
	LAYER VIA5 ;
		RECT -0.037500 -0.022500 0.037500 0.115 ;
	LAYER M6 ;
		RECT -0.037500 -0.097500 0.037500 0.375 ;
END VIA56_2cut_P2_SLN

VIA VIA56_2cut_P2_SLS DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M5 ;
		RECT -0.082500 -0.187500 0.082500 0.025 ;
	LAYER VIA5 ;
		RECT -0.037500 -0.172500 0.037500 0.015 ;
	LAYER M6 ;
		RECT -0.037500 -0.562500 0.037500 0.065 ;
END VIA56_2cut_P2_SLS

VIA VIA56_2cut_P3_N DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M5 ;
		RECT -0.082500 -0.037500 0.082500 0.125 ;
	LAYER VIA5 ;
		RECT -0.037500 -0.022500 0.037500 0.115 ;
	LAYER M6 ;
		RECT -0.037500 -0.082500 0.037500 0.155 ;
END VIA56_2cut_P3_N

VIA VIA56_2cut_P3_S DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M5 ;
		RECT -0.082500 -0.187500 0.082500 0.025 ;
	LAYER VIA5 ;
		RECT -0.037500 -0.172500 0.037500 0.015 ;
	LAYER M6 ;
		RECT -0.037500 -0.232500 0.037500 0.055 ;
END VIA56_2cut_P3_S

VIA VIA56_4cut DEFAULT
	RESISTANCE 3.000000 ;
	LAYER M5 ;
		RECT -0.180000 -0.135000 0.180000 0.09 ;
	LAYER VIA5 ;
		RECT -0.135000 -0.135000 -0.060000 -0.04 ;
		RECT 0.060000 -0.135000 0.135000 -0.04 ;
		RECT -0.135000 0.060000 -0.060000 0.09 ;
		RECT 0.060000 0.060000 0.135000 0.09 ;
	LAYER M6 ;
		RECT -0.135000 -0.180000 0.135000 0.12 ;
END VIA56_4cut

VIA VIA56_FBD_XEN DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M5 ;
		RECT -0.037500 -0.037500 0.247500 0.085 ;
	LAYER VIA5 ;
		RECT 0.007500 0.007500 0.202500 0.055 ;
	LAYER M6 ;
		RECT -0.037500 -0.037500 0.247500 0.085 ;
END VIA56_FBD_XEN

VIA VIA56_FBD_XES DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M5 ;
		RECT -0.037500 -0.127500 0.247500 0.025 ;
	LAYER VIA5 ;
		RECT 0.007500 -0.082500 0.202500 -0.005 ;
	LAYER M6 ;
		RECT -0.037500 -0.127500 0.247500 0.025 ;
END VIA56_FBD_XES

VIA VIA56_FBD_XWN DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M5 ;
		RECT -0.247500 -0.037500 0.037500 0.085 ;
	LAYER VIA5 ;
		RECT -0.202500 0.007500 -0.007500 0.055 ;
	LAYER M6 ;
		RECT -0.247500 -0.037500 0.037500 0.085 ;
END VIA56_FBD_XWN

VIA VIA56_FBD_XWS DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M5 ;
		RECT -0.247500 -0.127500 0.037500 0.025 ;
	LAYER VIA5 ;
		RECT -0.202500 -0.082500 -0.007500 -0.005 ;
	LAYER M6 ;
		RECT -0.247500 -0.127500 0.037500 0.025 ;
END VIA56_FBD_XWS

VIA VIA56_FBD_YEN DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M5 ;
		RECT -0.037500 -0.037500 0.127500 0.165 ;
	LAYER VIA5 ;
		RECT 0.007500 0.007500 0.082500 0.135 ;
	LAYER M6 ;
		RECT -0.037500 -0.037500 0.127500 0.165 ;
END VIA56_FBD_YEN

VIA VIA56_FBD_YES DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M5 ;
		RECT -0.037500 -0.247500 0.127500 0.025 ;
	LAYER VIA5 ;
		RECT 0.007500 -0.202500 0.082500 -0.005 ;
	LAYER M6 ;
		RECT -0.037500 -0.247500 0.127500 0.025 ;
END VIA56_FBD_YES

VIA VIA56_FBD_YWN DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M5 ;
		RECT -0.127500 -0.037500 0.037500 0.165 ;
	LAYER VIA5 ;
		RECT -0.082500 0.007500 -0.007500 0.135 ;
	LAYER M6 ;
		RECT -0.127500 -0.037500 0.037500 0.165 ;
END VIA56_FBD_YWN

VIA VIA56_FBD_YWS DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M5 ;
		RECT -0.127500 -0.247500 0.037500 0.025 ;
	LAYER VIA5 ;
		RECT -0.082500 -0.202500 -0.007500 -0.005 ;
	LAYER M6 ;
		RECT -0.127500 -0.247500 0.037500 0.025 ;
END VIA56_FBD_YWS

VIA VIA56_FBS DEFAULT
	RESISTANCE 12.000000 ;
	LAYER M5 ;
		RECT -0.082500 -0.082500 0.082500 0.055 ;
	LAYER VIA5 ;
		RECT -0.037500 -0.037500 0.037500 0.025 ;
	LAYER M6 ;
		RECT -0.082500 -0.082500 0.082500 0.055 ;
END VIA56_FBS

VIA VIA56_FBS_EN DEFAULT
	RESISTANCE 12.000000 ;
	LAYER M5 ;
		RECT -0.037500 -0.037500 0.127500 0.085 ;
	LAYER VIA5 ;
		RECT 0.007500 0.007500 0.082500 0.055 ;
	LAYER M6 ;
		RECT -0.037500 -0.037500 0.127500 0.085 ;
END VIA56_FBS_EN

VIA VIA56_FBS_ES DEFAULT
	RESISTANCE 12.000000 ;
	LAYER M5 ;
		RECT -0.037500 -0.127500 0.127500 0.025 ;
	LAYER VIA5 ;
		RECT 0.007500 -0.082500 0.082500 -0.005 ;
	LAYER M6 ;
		RECT -0.037500 -0.127500 0.127500 0.025 ;
END VIA56_FBS_ES

VIA VIA56_FBS_WN DEFAULT
	RESISTANCE 12.000000 ;
	LAYER M5 ;
		RECT -0.127500 -0.037500 0.037500 0.085 ;
	LAYER VIA5 ;
		RECT -0.082500 0.007500 -0.007500 0.055 ;
	LAYER M6 ;
		RECT -0.127500 -0.037500 0.037500 0.085 ;
END VIA56_FBS_WN

VIA VIA56_FBS_WS DEFAULT
	RESISTANCE 12.000000 ;
	LAYER M5 ;
		RECT -0.127500 -0.127500 0.037500 0.025 ;
	LAYER VIA5 ;
		RECT -0.082500 -0.082500 -0.007500 -0.005 ;
	LAYER M6 ;
		RECT -0.127500 -0.127500 0.037500 0.025 ;
END VIA56_FBS_WS

VIA VIA56_PBD_E DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M5 ;
		RECT -0.052500 -0.037500 0.262500 0.025 ;
	LAYER VIA5 ;
		RECT 0.007500 -0.037500 0.202500 0.025 ;
	LAYER M6 ;
		RECT -0.037500 -0.082500 0.247500 0.055 ;
END VIA56_PBD_E

VIA VIA56_PBD_N DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M5 ;
		RECT -0.037500 -0.052500 0.037500 0.175 ;
	LAYER VIA5 ;
		RECT -0.037500 0.007500 0.037500 0.135 ;
	LAYER M6 ;
		RECT -0.082500 -0.037500 0.082500 0.165 ;
END VIA56_PBD_N

VIA VIA56_PBD_S DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M5 ;
		RECT -0.037500 -0.262500 0.037500 0.035 ;
	LAYER VIA5 ;
		RECT -0.037500 -0.202500 0.037500 -0.005 ;
	LAYER M6 ;
		RECT -0.082500 -0.247500 0.082500 0.025 ;
END VIA56_PBD_S

VIA VIA56_PBD_W DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M5 ;
		RECT -0.262500 -0.037500 0.052500 0.025 ;
	LAYER VIA5 ;
		RECT -0.202500 -0.037500 -0.007500 0.025 ;
	LAYER M6 ;
		RECT -0.247500 -0.082500 0.037500 0.055 ;
END VIA56_PBD_W

VIA VIA56_PBS_H DEFAULT
	RESISTANCE 12.000000 ;
	LAYER M5 ;
		RECT -0.082500 -0.037500 0.082500 0.025 ;
	LAYER VIA5 ;
		RECT -0.037500 -0.037500 0.037500 0.025 ;
	LAYER M6 ;
		RECT -0.082500 -0.082500 0.082500 0.055 ;
END VIA56_PBS_H

VIA VIA56_PBS_V DEFAULT
	RESISTANCE 12.000000 ;
	LAYER M5 ;
		RECT -0.037500 -0.082500 0.037500 0.055 ;
	LAYER VIA5 ;
		RECT -0.037500 -0.037500 0.037500 0.025 ;
	LAYER M6 ;
		RECT -0.082500 -0.082500 0.082500 0.055 ;
END VIA56_PBS_V

VIA VIA56_FBD20_XEN DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M5 ;
		RECT -0.037500 -0.037500 0.217500 0.065 ;
	LAYER VIA5 ;
		RECT -0.007500 -0.007500 0.187500 0.045 ;
	LAYER M6 ;
		RECT -0.037500 -0.037500 0.217500 0.065 ;
END VIA56_FBD20_XEN

VIA VIA56_FBD20_XES DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M5 ;
		RECT -0.037500 -0.097500 0.217500 0.025 ;
	LAYER VIA5 ;
		RECT -0.007500 -0.067500 0.187500 0.005 ;
	LAYER M6 ;
		RECT -0.037500 -0.097500 0.217500 0.025 ;
END VIA56_FBD20_XES

VIA VIA56_FBD20_XWN DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M5 ;
		RECT -0.217500 -0.037500 0.037500 0.065 ;
	LAYER VIA5 ;
		RECT -0.187500 -0.007500 0.007500 0.045 ;
	LAYER M6 ;
		RECT -0.217500 -0.037500 0.037500 0.065 ;
END VIA56_FBD20_XWN

VIA VIA56_FBD20_XWS DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M5 ;
		RECT -0.217500 -0.097500 0.037500 0.025 ;
	LAYER VIA5 ;
		RECT -0.187500 -0.067500 0.007500 0.005 ;
	LAYER M6 ;
		RECT -0.217500 -0.097500 0.037500 0.025 ;
END VIA56_FBD20_XWS

VIA VIA56_FBD20_YEN DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M5 ;
		RECT -0.037500 -0.037500 0.097500 0.145 ;
	LAYER VIA5 ;
		RECT -0.007500 -0.007500 0.067500 0.125 ;
	LAYER M6 ;
		RECT -0.037500 -0.037500 0.097500 0.145 ;
END VIA56_FBD20_YEN

VIA VIA56_FBD20_YES DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M5 ;
		RECT -0.037500 -0.217500 0.097500 0.025 ;
	LAYER VIA5 ;
		RECT -0.007500 -0.187500 0.067500 0.005 ;
	LAYER M6 ;
		RECT -0.037500 -0.217500 0.097500 0.025 ;
END VIA56_FBD20_YES

VIA VIA56_FBD20_YWN DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M5 ;
		RECT -0.097500 -0.037500 0.037500 0.145 ;
	LAYER VIA5 ;
		RECT -0.067500 -0.007500 0.007500 0.125 ;
	LAYER M6 ;
		RECT -0.097500 -0.037500 0.037500 0.145 ;
END VIA56_FBD20_YWN

VIA VIA56_FBD20_YWS DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M5 ;
		RECT -0.097500 -0.217500 0.037500 0.025 ;
	LAYER VIA5 ;
		RECT -0.067500 -0.187500 0.007500 0.005 ;
	LAYER M6 ;
		RECT -0.097500 -0.217500 0.037500 0.025 ;
END VIA56_FBD20_YWS

VIA VIA56_FBD30_XEN DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M5 ;
		RECT -0.037500 -0.037500 0.187500 0.085 ;
	LAYER VIA5 ;
		RECT -0.022500 0.007500 0.172500 0.055 ;
	LAYER M6 ;
		RECT -0.037500 -0.037500 0.187500 0.085 ;
END VIA56_FBD30_XEN

VIA VIA56_FBD30_XES DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M5 ;
		RECT -0.037500 -0.127500 0.187500 0.025 ;
	LAYER VIA5 ;
		RECT -0.022500 -0.082500 0.172500 -0.005 ;
	LAYER M6 ;
		RECT -0.037500 -0.127500 0.187500 0.025 ;
END VIA56_FBD30_XES

VIA VIA56_FBD30_XWN DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M5 ;
		RECT -0.187500 -0.037500 0.037500 0.085 ;
	LAYER VIA5 ;
		RECT -0.172500 0.007500 0.022500 0.055 ;
	LAYER M6 ;
		RECT -0.187500 -0.037500 0.037500 0.085 ;
END VIA56_FBD30_XWN

VIA VIA56_FBD30_XWS DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M5 ;
		RECT -0.187500 -0.127500 0.037500 0.025 ;
	LAYER VIA5 ;
		RECT -0.172500 -0.082500 0.022500 -0.005 ;
	LAYER M6 ;
		RECT -0.187500 -0.127500 0.037500 0.025 ;
END VIA56_FBD30_XWS

VIA VIA56_FBD30_YEN DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M5 ;
		RECT -0.037500 -0.037500 0.127500 0.125 ;
	LAYER VIA5 ;
		RECT 0.007500 -0.022500 0.082500 0.115 ;
	LAYER M6 ;
		RECT -0.037500 -0.037500 0.127500 0.125 ;
END VIA56_FBD30_YEN

VIA VIA56_FBD30_YES DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M5 ;
		RECT -0.037500 -0.187500 0.127500 0.025 ;
	LAYER VIA5 ;
		RECT 0.007500 -0.172500 0.082500 0.015 ;
	LAYER M6 ;
		RECT -0.037500 -0.187500 0.127500 0.025 ;
END VIA56_FBD30_YES

VIA VIA56_FBD30_YWN DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M5 ;
		RECT -0.127500 -0.037500 0.037500 0.125 ;
	LAYER VIA5 ;
		RECT -0.082500 -0.022500 -0.007500 0.115 ;
	LAYER M6 ;
		RECT -0.127500 -0.037500 0.037500 0.125 ;
END VIA56_FBD30_YWN

VIA VIA56_FBD30_YWS DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M5 ;
		RECT -0.127500 -0.187500 0.037500 0.025 ;
	LAYER VIA5 ;
		RECT -0.082500 -0.172500 -0.007500 0.015 ;
	LAYER M6 ;
		RECT -0.127500 -0.187500 0.037500 0.025 ;
END VIA56_FBD30_YWS

VIA VIA56_PBDB_E DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M5 ;
		RECT -0.007500 -0.067500 0.247500 0.045 ;
	LAYER VIA5 ;
		RECT 0.022500 -0.037500 0.217500 0.025 ;
	LAYER M6 ;
		RECT -0.037500 -0.037500 0.277500 0.025 ;
END VIA56_PBDB_E

VIA VIA56_PBDB_N DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M5 ;
		RECT -0.067500 -0.007500 0.067500 0.165 ;
	LAYER VIA5 ;
		RECT -0.037500 0.022500 0.037500 0.145 ;
	LAYER M6 ;
		RECT -0.037500 -0.037500 0.037500 0.185 ;
END VIA56_PBDB_N

VIA VIA56_PBDB_S DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M5 ;
		RECT -0.067500 -0.247500 0.067500 0.005 ;
	LAYER VIA5 ;
		RECT -0.037500 -0.217500 0.037500 -0.015 ;
	LAYER M6 ;
		RECT -0.037500 -0.277500 0.037500 0.025 ;
END VIA56_PBDB_S

VIA VIA56_PBDB_W DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M5 ;
		RECT -0.247500 -0.067500 0.007500 0.045 ;
	LAYER VIA5 ;
		RECT -0.217500 -0.037500 -0.022500 0.025 ;
	LAYER M6 ;
		RECT -0.277500 -0.037500 0.037500 0.025 ;
END VIA56_PBDB_W

VIA VIA56_PBDU_E DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M5 ;
		RECT -0.067500 -0.037500 0.247500 0.025 ;
	LAYER VIA5 ;
		RECT -0.007500 -0.037500 0.187500 0.025 ;
	LAYER M6 ;
		RECT -0.037500 -0.067500 0.217500 0.045 ;
END VIA56_PBDU_E

VIA VIA56_PBDU_N DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M5 ;
		RECT -0.037500 -0.067500 0.037500 0.165 ;
	LAYER VIA5 ;
		RECT -0.037500 -0.007500 0.037500 0.125 ;
	LAYER M6 ;
		RECT -0.067500 -0.037500 0.067500 0.145 ;
END VIA56_PBDU_N

VIA VIA56_PBDU_S DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M5 ;
		RECT -0.037500 -0.247500 0.037500 0.045 ;
	LAYER VIA5 ;
		RECT -0.037500 -0.187500 0.037500 0.005 ;
	LAYER M6 ;
		RECT -0.067500 -0.217500 0.067500 0.025 ;
END VIA56_PBDU_S

VIA VIA56_PBDU_W DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M5 ;
		RECT -0.247500 -0.037500 0.067500 0.025 ;
	LAYER VIA5 ;
		RECT -0.187500 -0.037500 0.007500 0.025 ;
	LAYER M6 ;
		RECT -0.217500 -0.067500 0.037500 0.045 ;
END VIA56_PBDU_W

VIA VIA56_PBDE_E DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M5 ;
		RECT -0.037500 -0.037500 0.277500 0.025 ;
	LAYER VIA5 ;
		RECT 0.022500 -0.037500 0.217500 0.025 ;
	LAYER M6 ;
		RECT -0.037500 -0.037500 0.277500 0.025 ;
END VIA56_PBDE_E

VIA VIA56_PBDE_N DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M5 ;
		RECT -0.037500 -0.037500 0.037500 0.185 ;
	LAYER VIA5 ;
		RECT -0.037500 0.022500 0.037500 0.145 ;
	LAYER M6 ;
		RECT -0.037500 -0.037500 0.037500 0.185 ;
END VIA56_PBDE_N

VIA VIA56_PBDE_S DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M5 ;
		RECT -0.037500 -0.277500 0.037500 0.025 ;
	LAYER VIA5 ;
		RECT -0.037500 -0.217500 0.037500 -0.015 ;
	LAYER M6 ;
		RECT -0.037500 -0.277500 0.037500 0.025 ;
END VIA56_PBDE_S

VIA VIA56_PBDE_W DEFAULT
	RESISTANCE 6.750000 ;
	LAYER M5 ;
		RECT -0.277500 -0.037500 0.037500 0.025 ;
	LAYER VIA5 ;
		RECT -0.217500 -0.037500 -0.022500 0.025 ;
	LAYER M6 ;
		RECT -0.277500 -0.037500 0.037500 0.025 ;
END VIA56_PBDE_W

VIA VIA56_FBS25 DEFAULT
	RESISTANCE 12.000000 ;
	LAYER M5 ;
		RECT -0.075000 -0.075000 0.075000 0.05 ;
	LAYER VIA5 ;
		RECT -0.037500 -0.037500 0.037500 0.025 ;
	LAYER M6 ;
		RECT -0.075000 -0.075000 0.075000 0.05 ;
END VIA56_FBS25

VIA VIA56_FBS25_EN DEFAULT
	RESISTANCE 12.000000 ;
	LAYER M5 ;
		RECT -0.037500 -0.037500 0.112500 0.075 ;
	LAYER VIA5 ;
		RECT 0.000000 0.000000 0.075000 0.05 ;
	LAYER M6 ;
		RECT -0.037500 -0.037500 0.112500 0.075 ;
END VIA56_FBS25_EN

VIA VIA56_FBS25_ES DEFAULT
	RESISTANCE 12.000000 ;
	LAYER M5 ;
		RECT -0.037500 -0.112500 0.112500 0.025 ;
	LAYER VIA5 ;
		RECT 0.000000 -0.075000 0.075000 0 ;
	LAYER M6 ;
		RECT -0.037500 -0.112500 0.112500 0.025 ;
END VIA56_FBS25_ES

VIA VIA56_FBS25_WN DEFAULT
	RESISTANCE 12.000000 ;
	LAYER M5 ;
		RECT -0.112500 -0.037500 0.037500 0.075 ;
	LAYER VIA5 ;
		RECT -0.075000 0.000000 0.000000 0.05 ;
	LAYER M6 ;
		RECT -0.112500 -0.037500 0.037500 0.075 ;
END VIA56_FBS25_WN

VIA VIA56_FBS25_WS DEFAULT
	RESISTANCE 12.000000 ;
	LAYER M5 ;
		RECT -0.112500 -0.112500 0.037500 0.025 ;
	LAYER VIA5 ;
		RECT -0.075000 -0.075000 0.000000 0 ;
	LAYER M6 ;
		RECT -0.112500 -0.112500 0.037500 0.025 ;
END VIA56_FBS25_WS

VIA VIA56_PBSU_H DEFAULT
	RESISTANCE 12.000000 ;
	LAYER M5 ;
		RECT -0.082500 -0.037500 0.082500 0.025 ;
	LAYER VIA5 ;
		RECT -0.037500 -0.037500 0.037500 0.025 ;
	LAYER M6 ;
		RECT -0.052500 -0.075000 0.052500 0.05 ;
END VIA56_PBSU_H

VIA VIA56_PBSU_V DEFAULT
	RESISTANCE 12.000000 ;
	LAYER M5 ;
		RECT -0.037500 -0.082500 0.037500 0.055 ;
	LAYER VIA5 ;
		RECT -0.037500 -0.037500 0.037500 0.025 ;
	LAYER M6 ;
		RECT -0.075000 -0.052500 0.075000 0.035 ;
END VIA56_PBSU_V

VIA VIA56_PBSB_H DEFAULT
	RESISTANCE 12.000000 ;
	LAYER M5 ;
		RECT -0.075000 -0.052500 0.075000 0.035 ;
	LAYER VIA5 ;
		RECT -0.037500 -0.037500 0.037500 0.025 ;
	LAYER M6 ;
		RECT -0.037500 -0.082500 0.037500 0.055 ;
END VIA56_PBSB_H

VIA VIA56_PBSB_V DEFAULT
	RESISTANCE 12.000000 ;
	LAYER M5 ;
		RECT -0.052500 -0.075000 0.052500 0.05 ;
	LAYER VIA5 ;
		RECT -0.037500 -0.037500 0.037500 0.025 ;
	LAYER M6 ;
		RECT -0.082500 -0.037500 0.082500 0.025 ;
END VIA56_PBSB_V


VIA VIA67_1cut DEFAULT
	RESISTANCE 0.405000 ;
	LAYER M6 ;
		RECT -0.300000 -0.390000 0.300000 0.26 ;
	LAYER VIA6 ;
		RECT -0.270000 -0.270000 0.270000 0.18 ;
	LAYER M7 ;
		RECT -0.390000 -0.300000 0.390000 0.2 ;
END VIA67_1cut

VIA VIA67_1cut_H DEFAULT
	RESISTANCE 0.405000 ;
	LAYER M6 ;
		RECT -0.390000 -0.300000 0.390000 0.2 ;
	LAYER VIA6 ;
		RECT -0.270000 -0.270000 0.270000 0.18 ;
	LAYER M7 ;
		RECT -0.390000 -0.300000 0.390000 0.2 ;
END VIA67_1cut_H

VIA VIA67_1cut_V DEFAULT
	RESISTANCE 0.405000 ;
	LAYER M6 ;
		RECT -0.300000 -0.390000 0.300000 0.26 ;
	LAYER VIA6 ;
		RECT -0.270000 -0.270000 0.270000 0.18 ;
	LAYER M7 ;
		RECT -0.300000 -0.390000 0.300000 0.26 ;
END VIA67_1cut_V

VIA VIA67_2cut_P3_E DEFAULT
	RESISTANCE 0.202500 ;
	LAYER M6 ;
		RECT -0.300000 -0.390000 1.350000 0.26 ;
	LAYER VIA6 ;
		RECT -0.270000 -0.270000 0.270000 0.18 ;
		RECT 0.780000 -0.270000 1.320000 0.18 ;
	LAYER M7 ;
		RECT -0.390000 -0.300000 1.440000 0.2 ;
END VIA67_2cut_P3_E

VIA VIA67_2cut_P3_W DEFAULT
	RESISTANCE 0.202500 ;
	LAYER M6 ;
		RECT -1.350000 -0.390000 0.300000 0.26 ;
	LAYER VIA6 ;
		RECT -1.320000 -0.270000 -0.780000 0.18 ;
		RECT -0.270000 -0.270000 0.270000 0.18 ;
	LAYER M7 ;
		RECT -1.440000 -0.300000 0.390000 0.2 ;
END VIA67_2cut_P3_W

VIA VIA67_2cut_P1_N DEFAULT
	RESISTANCE 0.202500 ;
	LAYER M6 ;
		RECT -0.300000 -0.390000 0.300000 0.96 ;
	LAYER VIA6 ;
		RECT -0.270000 -0.270000 0.270000 0.18 ;
		RECT -0.270000 0.780000 0.270000 0.88 ;
	LAYER M7 ;
		RECT -0.390000 -0.300000 0.390000 0.9 ;
END VIA67_2cut_P1_N

VIA VIA67_2cut_P1_S DEFAULT
	RESISTANCE 0.202500 ;
	LAYER M6 ;
		RECT -0.300000 -1.440000 0.300000 0.26 ;
	LAYER VIA6 ;
		RECT -0.270000 -1.320000 0.270000 -0.52 ;
		RECT -0.270000 -0.270000 0.270000 0.18 ;
	LAYER M7 ;
		RECT -0.390000 -1.350000 0.390000 0.2 ;
END VIA67_2cut_P1_S

VIA VIA67_4cut DEFAULT
	RESISTANCE 0.101250 ;
	LAYER M6 ;
		RECT -0.975000 -1.065000 0.975000 0.71 ;
	LAYER VIA6 ;
		RECT -0.945000 -0.945000 -0.405000 -0.27 ;
		RECT 0.405000 -0.945000 0.945000 -0.27 ;
		RECT -0.945000 0.405000 -0.405000 0.63 ;
		RECT 0.405000 0.405000 0.945000 0.63 ;
	LAYER M7 ;
		RECT -1.065000 -0.975000 1.065000 0.65 ;
END VIA67_4cut

VIA VIA67_FBS DEFAULT
	RESISTANCE 0.405000 ;
	LAYER M6 ;
		RECT -0.390000 -0.390000 0.390000 0.26 ;
	LAYER VIA6 ;
		RECT -0.270000 -0.270000 0.270000 0.18 ;
	LAYER M7 ;
		RECT -0.390000 -0.390000 0.390000 0.26 ;
END VIA67_FBS


VIA VIA78_1cut DEFAULT
	RESISTANCE 0.405000 ;
	LAYER M7 ;
		RECT -0.390000 -0.390000 0.390000 0.26 ;
	LAYER VIA7 ;
		RECT -0.270000 -0.270000 0.270000 0.18 ;
	LAYER M8 ;
		RECT -1.500000 -1.500000 1.500000 1 ;
END VIA78_1cut

VIA VIA78_2cut_P1_E DEFAULT
	RESISTANCE 0.202500 ;
	LAYER M7 ;
		RECT -0.390000 -0.390000 1.440000 0.26 ;
	LAYER VIA7 ;
		RECT -0.270000 -0.270000 0.270000 0.18 ;
		RECT 0.780000 -0.270000 1.320000 0.18 ;
	LAYER M8 ;
		RECT -0.975000 -1.500000 2.025000 1 ;
END VIA78_2cut_P1_E

VIA VIA78_2cut_P1_W DEFAULT
	RESISTANCE 0.202500 ;
	LAYER M7 ;
		RECT -1.440000 -0.390000 0.390000 0.26 ;
	LAYER VIA7 ;
		RECT -1.320000 -0.270000 -0.780000 0.18 ;
		RECT -0.270000 -0.270000 0.270000 0.18 ;
	LAYER M8 ;
		RECT -2.025000 -1.500000 0.975000 1 ;
END VIA78_2cut_P1_W

VIA VIA78_2cut_P1_N DEFAULT
	RESISTANCE 0.202500 ;
	LAYER M7 ;
		RECT -0.390000 -0.390000 0.390000 0.96 ;
	LAYER VIA7 ;
		RECT -0.270000 -0.270000 0.270000 0.18 ;
		RECT -0.270000 0.780000 0.270000 0.88 ;
	LAYER M8 ;
		RECT -1.500000 -0.975000 1.500000 1.35 ;
END VIA78_2cut_P1_N

VIA VIA78_2cut_P1_S DEFAULT
	RESISTANCE 0.202500 ;
	LAYER M7 ;
		RECT -0.390000 -1.440000 0.390000 0.26 ;
	LAYER VIA7 ;
		RECT -0.270000 -1.320000 0.270000 -0.52 ;
		RECT -0.270000 -0.270000 0.270000 0.18 ;
	LAYER M8 ;
		RECT -1.500000 -2.025000 1.500000 0.65 ;
END VIA78_2cut_P1_S


VIA VIA8AP_1cut DEFAULT
	RESISTANCE 0.096000 ;
	LAYER M8 ;
		RECT -3.000000 -3.000000 3.000000 2 ;
	LAYER RV ;
		RECT -2.250000 -2.250000 2.250000 1.5 ;
	LAYER AP ;
		RECT -3.000000 -3.000000 3.000000 2 ;
END VIA8AP_1cut


VIARULE VIAGEN12 GENERATE
    LAYER M1 ;
        ENCLOSURE 0.045000 0.000000 ;
        WIDTH 0.075000 TO 6.750000 ;
    LAYER M2 ;
        ENCLOSURE 0.045000 0.000000 ;
        WIDTH 0.075000 TO 6.750000 ;
    LAYER VIA1 ;
		RECT -0.037500 -0.037500 0.037500 0.025 ;
        SPACING 0.195000 BY 0.195000 ;
END VIAGEN12


VIARULE VIAGEN12_RECT GENERATE
    LAYER M1 ;
        ENCLOSURE 0.060000 0.000000 ;
        WIDTH 0.075000 TO 6.750000 ;
    LAYER M2 ;
        ENCLOSURE 0.060000 0.000000 ;
        WIDTH 0.075000 TO 6.750000 ;
    LAYER VIA1 ;
		RECT -0.037500 -0.037500 0.157500 0.025000 ;
        SPACING 0.315000 BY 0.195000 ;
END VIAGEN12_RECT


VIARULE VIAGEN23 GENERATE
    LAYER M2 ;
        ENCLOSURE 0.045000 0.000000 ;
        WIDTH 0.075000 TO 6.750000 ;
    LAYER M3 ;
        ENCLOSURE 0.045000 0.000000 ;
        WIDTH 0.075000 TO 6.750000 ;
    LAYER VIA2 ;
		RECT -0.037500 -0.037500 0.037500 0.025 ;
        SPACING 0.195000 BY 0.195000 ;
END VIAGEN23


VIARULE VIAGEN23_RECT GENERATE
    LAYER M2 ;
        ENCLOSURE 0.060000 0.000000 ;
        WIDTH 0.075000 TO 6.750000 ;
    LAYER M3 ;
        ENCLOSURE 0.060000 0.000000 ;
        WIDTH 0.075000 TO 6.750000 ;
    LAYER VIA2 ;
		RECT -0.037500 -0.037500 0.157500 0.025000 ;
        SPACING 0.315000 BY 0.195000 ;
END VIAGEN23_RECT


VIARULE VIAGEN34 GENERATE
    LAYER M3 ;
        ENCLOSURE 0.045000 0.000000 ;
        WIDTH 0.075000 TO 6.750000 ;
    LAYER M4 ;
        ENCLOSURE 0.045000 0.000000 ;
        WIDTH 0.075000 TO 6.750000 ;
    LAYER VIA3 ;
		RECT -0.037500 -0.037500 0.037500 0.025 ;
        SPACING 0.195000 BY 0.195000 ;
END VIAGEN34


VIARULE VIAGEN34_RECT GENERATE
    LAYER M3 ;
        ENCLOSURE 0.060000 0.000000 ;
        WIDTH 0.075000 TO 6.750000 ;
    LAYER M4 ;
        ENCLOSURE 0.060000 0.000000 ;
        WIDTH 0.075000 TO 6.750000 ;
    LAYER VIA3 ;
		RECT -0.037500 -0.037500 0.157500 0.025000 ;
        SPACING 0.315000 BY 0.195000 ;
END VIAGEN34_RECT


VIARULE VIAGEN45 GENERATE
    LAYER M4 ;
        ENCLOSURE 0.045000 0.000000 ;
        WIDTH 0.075000 TO 6.750000 ;
    LAYER M5 ;
        ENCLOSURE 0.045000 0.000000 ;
        WIDTH 0.075000 TO 6.750000 ;
    LAYER VIA4 ;
		RECT -0.037500 -0.037500 0.037500 0.025 ;
        SPACING 0.195000 BY 0.195000 ;
END VIAGEN45


VIARULE VIAGEN45_RECT GENERATE
    LAYER M4 ;
        ENCLOSURE 0.060000 0.000000 ;
        WIDTH 0.075000 TO 6.750000 ;
    LAYER M5 ;
        ENCLOSURE 0.060000 0.000000 ;
        WIDTH 0.075000 TO 6.750000 ;
    LAYER VIA4 ;
		RECT -0.037500 -0.037500 0.157500 0.025000 ;
        SPACING 0.315000 BY 0.195000 ;
END VIAGEN45_RECT


VIARULE VIAGEN56 GENERATE
    LAYER M5 ;
        ENCLOSURE 0.045000 0.000000 ;
        WIDTH 0.075000 TO 6.750000 ;
    LAYER M6 ;
        ENCLOSURE 0.045000 0.000000 ;
        WIDTH 0.075000 TO 6.750000 ;
    LAYER VIA5 ;
		RECT -0.037500 -0.037500 0.037500 0.025 ;
        SPACING 0.195000 BY 0.195000 ;
END VIAGEN56


VIARULE VIAGEN56_RECT GENERATE
    LAYER M5 ;
        ENCLOSURE 0.060000 0.000000 ;
        WIDTH 0.075000 TO 6.750000 ;
    LAYER M6 ;
        ENCLOSURE 0.060000 0.000000 ;
        WIDTH 0.075000 TO 6.750000 ;
    LAYER VIA5 ;
		RECT -0.037500 -0.037500 0.157500 0.025000 ;
        SPACING 0.315000 BY 0.195000 ;
END VIAGEN56_RECT


VIARULE VIAGEN67 GENERATE
    LAYER M6 ;
        ENCLOSURE 0.120000 0.030000 ;
        WIDTH 0.075000 TO 6.750000 ;
    LAYER M7 ;
        ENCLOSURE 0.120000 0.030000 ;
        WIDTH 0.600000 TO 18.000000 ;
    LAYER VIA6 ;
		RECT -0.270000 -0.270000 0.270000 0.18 ;
        SPACING 1.350000 BY 1.350000 ;
END VIAGEN67


VIARULE VIAGEN78 GENERATE
    LAYER M7 ;
        ENCLOSURE 0.120000 0.120000 ;
        WIDTH 0.600000 TO 18.000000 ;
    LAYER M8 ;
        ENCLOSURE 0.120000 0.120000 ;
        WIDTH 3.000000 TO 18.000000 ;
    LAYER VIA7 ;
		RECT -0.270000 -0.270000 0.270000 0.18 ;
        SPACING 1.350000 BY 1.350000 ;
END VIAGEN78


VIARULE VIAGEN8AP GENERATE
    LAYER M8 ;
        ENCLOSURE 0.750000 0.750000 ;
        WIDTH 3.000000 TO 18.000000 ;
    LAYER AP ;
        ENCLOSURE 0.750000 0.750000 ;
        WIDTH 3.000000 TO 52.500000 ;
    LAYER RV ;
		RECT -2.250000 -2.250000 2.250000 1.500000 ;
        SPACING 7.500000 BY 7.500000 ;
END VIAGEN8AP

MACRO AN2_0010
    CLASS CORE ;
    FOREIGN AN2_0010 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.2000 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 3.4125 0.2775 3.5700 0.3975 ;
        RECT 3.4125 0.6525 3.5700 0.7725 ;
        RECT 3.0975 0.2775 3.4125 0.7725 ;
        RECT 2.9400 0.2775 3.0975 0.3975 ;
        RECT 2.9400 0.6525 3.0975 0.7725 ;
        VIA 3.4125 0.3375 VIA12_slot ;
        VIA 3.4125 0.7125 VIA12_slot ;
        VIA 3.0975 0.3375 VIA12_slot ;
        VIA 3.0975 0.7125 VIA12_slot ;
        END
    END Z
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.3375 0.4125 1.3125 0.5325 ;
        RECT 0.1725 0.4125 0.3375 0.6375 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.8000 0.4350 1.9050 0.6375 ;
        RECT 1.3050 0.5625 1.8000 0.6375 ;
        VIA 1.8525 0.5400 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 4.1550 -0.0750 4.2000 0.0750 ;
        RECT 4.0350 -0.0750 4.1550 0.2925 ;
        RECT 3.7350 -0.0750 4.0350 0.0750 ;
        RECT 3.6150 -0.0750 3.7350 0.2025 ;
        RECT 3.3150 -0.0750 3.6150 0.0750 ;
        RECT 3.1950 -0.0750 3.3150 0.2025 ;
        RECT 2.8950 -0.0750 3.1950 0.0750 ;
        RECT 2.7750 -0.0750 2.8950 0.2025 ;
        RECT 2.4675 -0.0750 2.7750 0.0750 ;
        RECT 2.3625 -0.0750 2.4675 0.2400 ;
        RECT 1.2150 -0.0750 2.3625 0.0750 ;
        RECT 1.0950 -0.0750 1.2150 0.1875 ;
        RECT 0.7950 -0.0750 1.0950 0.0750 ;
        RECT 0.6750 -0.0750 0.7950 0.1875 ;
        RECT 0.3750 -0.0750 0.6750 0.0750 ;
        RECT 0.2550 -0.0750 0.3750 0.1875 ;
        RECT 0.0000 -0.0750 0.2550 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 4.1550 0.9750 4.2000 1.1250 ;
        RECT 4.0350 0.6600 4.1550 1.1250 ;
        RECT 3.7350 0.9750 4.0350 1.1250 ;
        RECT 3.6150 0.8475 3.7350 1.1250 ;
        RECT 3.3150 0.9750 3.6150 1.1250 ;
        RECT 3.1950 0.8475 3.3150 1.1250 ;
        RECT 2.8950 0.9750 3.1950 1.1250 ;
        RECT 2.7750 0.8475 2.8950 1.1250 ;
        RECT 2.4750 0.9750 2.7750 1.1250 ;
        RECT 2.3550 0.8175 2.4750 1.1250 ;
        RECT 2.2650 0.9750 2.3550 1.1250 ;
        RECT 2.1450 0.8175 2.2650 1.1250 ;
        RECT 1.8375 0.9750 2.1450 1.1250 ;
        RECT 1.7325 0.8250 1.8375 1.1250 ;
        RECT 1.4175 0.9750 1.7325 1.1250 ;
        RECT 1.3125 0.8250 1.4175 1.1250 ;
        RECT 0.9975 0.9750 1.3125 1.1250 ;
        RECT 0.8925 0.8250 0.9975 1.1250 ;
        RECT 0.5850 0.9750 0.8925 1.1250 ;
        RECT 0.4650 0.8625 0.5850 1.1250 ;
        RECT 0.1425 0.9750 0.4650 1.1250 ;
        RECT 0.0675 0.7800 0.1425 1.1250 ;
        RECT 0.0000 0.9750 0.0675 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 4.0650 0.2175 4.1250 0.2775 ;
        RECT 4.0650 0.6675 4.1250 0.7275 ;
        RECT 4.0650 0.8325 4.1250 0.8925 ;
        RECT 3.9600 0.4800 4.0200 0.5400 ;
        RECT 3.8550 0.3075 3.9150 0.3675 ;
        RECT 3.8550 0.6825 3.9150 0.7425 ;
        RECT 3.7500 0.4800 3.8100 0.5400 ;
        RECT 3.6450 0.1350 3.7050 0.1950 ;
        RECT 3.6450 0.8550 3.7050 0.9150 ;
        RECT 3.5400 0.4800 3.6000 0.5400 ;
        RECT 3.4350 0.3075 3.4950 0.3675 ;
        RECT 3.4350 0.6825 3.4950 0.7425 ;
        RECT 3.3300 0.4800 3.3900 0.5400 ;
        RECT 3.2250 0.1350 3.2850 0.1950 ;
        RECT 3.2250 0.8550 3.2850 0.9150 ;
        RECT 3.1200 0.4800 3.1800 0.5400 ;
        RECT 3.0150 0.3075 3.0750 0.3675 ;
        RECT 3.0150 0.6825 3.0750 0.7425 ;
        RECT 2.9100 0.4800 2.9700 0.5400 ;
        RECT 2.8050 0.1350 2.8650 0.1950 ;
        RECT 2.8050 0.8550 2.8650 0.9150 ;
        RECT 2.7000 0.4800 2.7600 0.5400 ;
        RECT 2.5950 0.3075 2.6550 0.3675 ;
        RECT 2.5950 0.6825 2.6550 0.7425 ;
        RECT 2.4900 0.4800 2.5500 0.5400 ;
        RECT 2.3850 0.1575 2.4450 0.2175 ;
        RECT 2.3850 0.8325 2.4450 0.8925 ;
        RECT 2.1750 0.1725 2.2350 0.2325 ;
        RECT 2.1750 0.8325 2.2350 0.8925 ;
        RECT 2.0700 0.4800 2.1300 0.5400 ;
        RECT 1.9650 0.3000 2.0250 0.3600 ;
        RECT 1.9650 0.7800 2.0250 0.8400 ;
        RECT 1.8600 0.4800 1.9200 0.5400 ;
        RECT 1.7550 0.1575 1.8150 0.2175 ;
        RECT 1.7550 0.8550 1.8150 0.9150 ;
        RECT 1.6500 0.4800 1.7100 0.5400 ;
        RECT 1.5450 0.3000 1.6050 0.3600 ;
        RECT 1.5450 0.6750 1.6050 0.7350 ;
        RECT 1.4400 0.4800 1.5000 0.5400 ;
        RECT 1.3350 0.1575 1.3950 0.2175 ;
        RECT 1.3350 0.8550 1.3950 0.9150 ;
        RECT 1.2225 0.4650 1.2825 0.5250 ;
        RECT 1.1250 0.1275 1.1850 0.1875 ;
        RECT 1.1250 0.6750 1.1850 0.7350 ;
        RECT 1.0200 0.4650 1.0800 0.5250 ;
        RECT 0.9150 0.2700 0.9750 0.3300 ;
        RECT 0.9150 0.8550 0.9750 0.9150 ;
        RECT 0.8100 0.4650 0.8700 0.5250 ;
        RECT 0.7050 0.1275 0.7650 0.1875 ;
        RECT 0.7050 0.8100 0.7650 0.8700 ;
        RECT 0.6000 0.4650 0.6600 0.5250 ;
        RECT 0.4950 0.2700 0.5550 0.3300 ;
        RECT 0.4950 0.8625 0.5550 0.9225 ;
        RECT 0.3900 0.4650 0.4500 0.5250 ;
        RECT 0.0750 0.8325 0.1350 0.8925 ;
        RECT 0.2850 0.1275 0.3450 0.1875 ;
        RECT 0.2850 0.8100 0.3450 0.8700 ;
        RECT 0.1800 0.4650 0.2400 0.5250 ;
        RECT 0.0750 0.2100 0.1350 0.2700 ;
        LAYER M1 ;
        RECT 2.4525 0.4725 4.0950 0.5475 ;
        RECT 2.5875 0.2775 3.9300 0.3975 ;
        RECT 2.5875 0.6525 3.9300 0.7725 ;
        RECT 2.3775 0.3300 2.4525 0.7425 ;
        RECT 2.0700 0.3300 2.3775 0.4050 ;
        RECT 2.0325 0.6675 2.3775 0.7425 ;
        RECT 2.1450 0.1500 2.2575 0.2550 ;
        RECT 1.4100 0.4800 2.2575 0.5850 ;
        RECT 1.3650 0.1500 2.1450 0.2250 ;
        RECT 1.5150 0.3000 2.0700 0.4050 ;
        RECT 1.9575 0.6675 2.0325 0.8700 ;
        RECT 0.7875 0.6675 1.9575 0.7425 ;
        RECT 1.2900 0.1500 1.3650 0.3375 ;
        RECT 0.1425 0.2625 1.2900 0.3375 ;
        RECT 0.6825 0.6675 0.7875 0.9000 ;
        RECT 0.3675 0.7125 0.6825 0.7875 ;
        RECT 0.2625 0.7125 0.3675 0.9000 ;
        RECT 0.0675 0.1800 0.1425 0.3375 ;
        LAYER M2 ;
        RECT 3.4425 0.2775 3.5700 0.3975 ;
        RECT 3.4425 0.6525 3.5700 0.7725 ;
        RECT 2.9400 0.2775 3.0675 0.3975 ;
        RECT 2.9400 0.6525 3.0675 0.7725 ;
    END
END AN2_0010


MACRO AN2_0011
    CLASS CORE ;
    FOREIGN AN2_0011 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.0500 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.9375 0.2925 1.0125 0.7425 ;
        RECT 0.6750 0.2925 0.9375 0.3675 ;
        RECT 0.7725 0.6675 0.9375 0.7425 ;
        RECT 0.6975 0.6675 0.7725 0.8550 ;
        END
    END Z
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.1875 0.2625 0.6525 0.3375 ;
        VIA 0.4800 0.3000 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.1875 0.4125 0.6525 0.4875 ;
        VIA 0.2700 0.4500 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.0050 -0.0750 1.0500 0.0750 ;
        RECT 0.8850 -0.0750 1.0050 0.2175 ;
        RECT 0.5925 -0.0750 0.8850 0.0750 ;
        RECT 0.4575 -0.0750 0.5925 0.1800 ;
        RECT 0.0000 -0.0750 0.4575 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.0050 0.9750 1.0500 1.1250 ;
        RECT 0.8850 0.8175 1.0050 1.1250 ;
        RECT 0.5850 0.9750 0.8850 1.1250 ;
        RECT 0.4650 0.8325 0.5850 1.1250 ;
        RECT 0.1650 0.9750 0.4650 1.1250 ;
        RECT 0.0450 0.8250 0.1650 1.1250 ;
        RECT 0.0000 0.9750 0.0450 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 0.9150 0.1575 0.9750 0.2175 ;
        RECT 0.9150 0.8325 0.9750 0.8925 ;
        RECT 0.8025 0.4950 0.8625 0.5550 ;
        RECT 0.7050 0.3000 0.7650 0.3600 ;
        RECT 0.7050 0.7650 0.7650 0.8250 ;
        RECT 0.6000 0.4950 0.6600 0.5550 ;
        RECT 0.4950 0.1200 0.5550 0.1800 ;
        RECT 0.4950 0.8550 0.5550 0.9150 ;
        RECT 0.3975 0.4800 0.4575 0.5400 ;
        RECT 0.2850 0.8175 0.3450 0.8775 ;
        RECT 0.1875 0.4800 0.2475 0.5400 ;
        RECT 0.0750 0.1575 0.1350 0.2175 ;
        RECT 0.0750 0.8325 0.1350 0.8925 ;
        LAYER M1 ;
        RECT 0.6225 0.4650 0.8625 0.5850 ;
        RECT 0.5475 0.4650 0.6225 0.7500 ;
        RECT 0.4725 0.2550 0.5625 0.3450 ;
        RECT 0.3675 0.6750 0.5475 0.7500 ;
        RECT 0.3975 0.2550 0.4725 0.5700 ;
        RECT 0.2625 0.6750 0.3675 0.9000 ;
        RECT 0.1875 0.3375 0.3225 0.6000 ;
        RECT 0.1125 0.6750 0.2625 0.7500 ;
        RECT 0.1125 0.1500 0.1650 0.2250 ;
        RECT 0.0375 0.1500 0.1125 0.7500 ;
    END
END AN2_0011


MACRO AN2_0100
    CLASS CORE ;
    FOREIGN AN2_0100 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.1500 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 2.3625 0.2625 2.5200 0.3825 ;
        RECT 2.3625 0.6600 2.5200 0.7800 ;
        RECT 2.0475 0.2625 2.3625 0.7800 ;
        RECT 1.8900 0.2625 2.0475 0.3825 ;
        RECT 1.8900 0.6600 2.0475 0.7800 ;
        VIA 2.3625 0.3225 VIA12_slot ;
        VIA 2.3625 0.7200 VIA12_slot ;
        VIA 2.0475 0.3225 VIA12_slot ;
        VIA 2.0475 0.7200 VIA12_slot ;
        END
    END Z
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.5700 0.4125 1.0350 0.4875 ;
        VIA 0.6750 0.4500 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.1275 0.5625 1.1250 0.6375 ;
        VIA 1.0425 0.6000 VIA12_square ;
        VIA 0.2100 0.6000 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 3.0825 -0.0750 3.1500 0.0750 ;
        RECT 3.0075 -0.0750 3.0825 0.2925 ;
        RECT 2.6850 -0.0750 3.0075 0.0750 ;
        RECT 2.5650 -0.0750 2.6850 0.1875 ;
        RECT 2.2650 -0.0750 2.5650 0.0750 ;
        RECT 2.1450 -0.0750 2.2650 0.1875 ;
        RECT 1.8450 -0.0750 2.1450 0.0750 ;
        RECT 1.7250 -0.0750 1.8450 0.1875 ;
        RECT 1.4175 -0.0750 1.7250 0.0750 ;
        RECT 1.3125 -0.0750 1.4175 0.2325 ;
        RECT 0.5625 -0.0750 1.3125 0.0750 ;
        RECT 0.4875 -0.0750 0.5625 0.2775 ;
        RECT 0.0000 -0.0750 0.4875 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 3.0825 0.9750 3.1500 1.1250 ;
        RECT 3.0075 0.6375 3.0825 1.1250 ;
        RECT 2.6850 0.9750 3.0075 1.1250 ;
        RECT 2.5650 0.8550 2.6850 1.1250 ;
        RECT 2.2650 0.9750 2.5650 1.1250 ;
        RECT 2.1450 0.8550 2.2650 1.1250 ;
        RECT 1.8450 0.9750 2.1450 1.1250 ;
        RECT 1.7250 0.8550 1.8450 1.1250 ;
        RECT 1.4250 0.9750 1.7250 1.1250 ;
        RECT 1.3050 0.8625 1.4250 1.1250 ;
        RECT 1.0050 0.9750 1.3050 1.1250 ;
        RECT 0.8850 0.8625 1.0050 1.1250 ;
        RECT 0.5850 0.9750 0.8850 1.1250 ;
        RECT 0.4650 0.8625 0.5850 1.1250 ;
        RECT 0.1575 0.9750 0.4650 1.1250 ;
        RECT 0.0525 0.8100 0.1575 1.1250 ;
        RECT 0.0000 0.9750 0.0525 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 3.0150 0.1875 3.0750 0.2475 ;
        RECT 3.0150 0.6675 3.0750 0.7275 ;
        RECT 3.0150 0.8325 3.0750 0.8925 ;
        RECT 2.9100 0.4650 2.9700 0.5250 ;
        RECT 2.8050 0.2850 2.8650 0.3450 ;
        RECT 2.8050 0.6900 2.8650 0.7500 ;
        RECT 2.7000 0.4650 2.7600 0.5250 ;
        RECT 2.5950 0.1275 2.6550 0.1875 ;
        RECT 2.5950 0.8625 2.6550 0.9225 ;
        RECT 2.4900 0.4650 2.5500 0.5250 ;
        RECT 2.3850 0.2850 2.4450 0.3450 ;
        RECT 2.3850 0.6900 2.4450 0.7500 ;
        RECT 2.2800 0.4650 2.3400 0.5250 ;
        RECT 2.1750 0.1275 2.2350 0.1875 ;
        RECT 2.1750 0.8625 2.2350 0.9225 ;
        RECT 2.0700 0.4650 2.1300 0.5250 ;
        RECT 1.9650 0.2850 2.0250 0.3450 ;
        RECT 1.9650 0.6900 2.0250 0.7500 ;
        RECT 1.8600 0.4650 1.9200 0.5250 ;
        RECT 1.7550 0.1275 1.8150 0.1875 ;
        RECT 1.7550 0.8625 1.8150 0.9225 ;
        RECT 1.6500 0.4650 1.7100 0.5250 ;
        RECT 1.5450 0.2850 1.6050 0.3450 ;
        RECT 1.5450 0.6900 1.6050 0.7500 ;
        RECT 1.4400 0.4650 1.5000 0.5250 ;
        RECT 1.3350 0.1500 1.3950 0.2100 ;
        RECT 1.3350 0.8700 1.3950 0.9300 ;
        RECT 1.2300 0.4800 1.2900 0.5400 ;
        RECT 1.1250 0.7200 1.1850 0.7800 ;
        RECT 1.0200 0.4875 1.0800 0.5475 ;
        RECT 0.9150 0.1575 0.9750 0.2175 ;
        RECT 0.9150 0.8700 0.9750 0.9300 ;
        RECT 0.8100 0.4875 0.8700 0.5475 ;
        RECT 0.7050 0.7200 0.7650 0.7800 ;
        RECT 0.6000 0.4800 0.6600 0.5400 ;
        RECT 0.4950 0.1875 0.5550 0.2475 ;
        RECT 0.4950 0.8700 0.5550 0.9300 ;
        RECT 0.3900 0.4800 0.4500 0.5400 ;
        RECT 0.2850 0.8175 0.3450 0.8775 ;
        RECT 0.1800 0.4800 0.2400 0.5400 ;
        RECT 0.0750 0.1875 0.1350 0.2475 ;
        RECT 0.0750 0.8325 0.1350 0.8925 ;
        LAYER M1 ;
        RECT 1.4625 0.4575 3.0000 0.5325 ;
        RECT 1.5225 0.2625 2.8875 0.3825 ;
        RECT 1.5375 0.6600 2.8875 0.7800 ;
        RECT 1.3875 0.4575 1.4625 0.7875 ;
        RECT 0.3675 0.7125 1.3875 0.7875 ;
        RECT 1.2300 0.3150 1.3050 0.5700 ;
        RECT 0.7125 0.3150 1.2300 0.3900 ;
        RECT 0.8025 0.1500 1.1925 0.2400 ;
        RECT 0.9600 0.4650 1.1250 0.6375 ;
        RECT 0.7875 0.4650 0.9600 0.5700 ;
        RECT 0.6375 0.3150 0.7125 0.5625 ;
        RECT 0.3675 0.4575 0.6375 0.5625 ;
        RECT 0.0675 0.1500 0.3825 0.2775 ;
        RECT 0.2625 0.7125 0.3675 0.9000 ;
        RECT 0.1275 0.4200 0.2925 0.6375 ;
        LAYER VIA1 ;
        RECT 1.3875 0.5025 1.4625 0.5775 ;
        RECT 1.0725 0.1650 1.1475 0.2400 ;
        RECT 0.2625 0.1650 0.3375 0.2400 ;
        LAYER M2 ;
        RECT 2.3925 0.2625 2.5200 0.3825 ;
        RECT 2.3925 0.6600 2.5200 0.7800 ;
        RECT 1.8900 0.2625 2.0175 0.3825 ;
        RECT 1.8900 0.6600 2.0175 0.7800 ;
        RECT 1.3725 0.2625 1.4775 0.6225 ;
        RECT 1.1925 0.2625 1.3725 0.3375 ;
        RECT 1.1175 0.1650 1.1925 0.3375 ;
        RECT 0.2175 0.1650 1.1175 0.2400 ;
    END
END AN2_0100


MACRO AN2_0111
    CLASS CORE ;
    FOREIGN AN2_0111 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.8900 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 1.2075 0.2625 1.5225 0.7500 ;
        VIA 1.3650 0.3450 VIA12_slot ;
        VIA 1.3650 0.6675 VIA12_slot ;
        END
    END Z
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.8100 0.3075 0.8850 0.5700 ;
        RECT 0.2925 0.3075 0.8100 0.3825 ;
        RECT 0.2175 0.3075 0.2925 0.5550 ;
        RECT 0.1425 0.4650 0.2175 0.5550 ;
        RECT 0.0675 0.4650 0.1425 0.6825 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.8175 0.7125 1.0575 0.7875 ;
        RECT 0.7425 0.5625 0.8175 0.7875 ;
        RECT 0.4275 0.5625 0.7425 0.6375 ;
        VIA 0.6225 0.6000 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.8225 -0.0750 1.8900 0.0750 ;
        RECT 1.7475 -0.0750 1.8225 0.3150 ;
        RECT 1.4250 -0.0750 1.7475 0.0750 ;
        RECT 1.3050 -0.0750 1.4250 0.2100 ;
        RECT 0.9975 -0.0750 1.3050 0.0750 ;
        RECT 0.8925 -0.0750 0.9975 0.2325 ;
        RECT 0.1425 -0.0750 0.8925 0.0750 ;
        RECT 0.0675 -0.0750 0.1425 0.2775 ;
        RECT 0.0000 -0.0750 0.0675 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.8225 0.9750 1.8900 1.1250 ;
        RECT 1.7475 0.6375 1.8225 1.1250 ;
        RECT 1.4025 0.9750 1.7475 1.1250 ;
        RECT 1.3275 0.8175 1.4025 1.1250 ;
        RECT 1.0050 0.9750 1.3275 1.1250 ;
        RECT 0.8850 0.8625 1.0050 1.1250 ;
        RECT 0.5850 0.9750 0.8850 1.1250 ;
        RECT 0.4650 0.8625 0.5850 1.1250 ;
        RECT 0.1575 0.9750 0.4650 1.1250 ;
        RECT 0.0525 0.8100 0.1575 1.1250 ;
        RECT 0.0000 0.9750 0.0525 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.7550 0.2250 1.8150 0.2850 ;
        RECT 1.7550 0.6675 1.8150 0.7275 ;
        RECT 1.7550 0.8325 1.8150 0.8925 ;
        RECT 1.6500 0.4650 1.7100 0.5250 ;
        RECT 1.5450 0.2250 1.6050 0.2850 ;
        RECT 1.5450 0.7200 1.6050 0.7800 ;
        RECT 1.4400 0.4650 1.5000 0.5250 ;
        RECT 1.3350 0.1275 1.3950 0.1875 ;
        RECT 1.3350 0.8475 1.3950 0.9075 ;
        RECT 1.2300 0.4650 1.2900 0.5250 ;
        RECT 1.1250 0.2250 1.1850 0.2850 ;
        RECT 1.1250 0.7200 1.1850 0.7800 ;
        RECT 1.0200 0.4650 1.0800 0.5250 ;
        RECT 0.9150 0.1500 0.9750 0.2100 ;
        RECT 0.9150 0.8700 0.9750 0.9300 ;
        RECT 0.8100 0.4800 0.8700 0.5400 ;
        RECT 0.7050 0.7200 0.7650 0.7800 ;
        RECT 0.6000 0.4800 0.6600 0.5400 ;
        RECT 0.4950 0.1575 0.5550 0.2175 ;
        RECT 0.4950 0.8700 0.5550 0.9300 ;
        RECT 0.3900 0.4800 0.4500 0.5400 ;
        RECT 0.2850 0.8175 0.3450 0.8775 ;
        RECT 0.1800 0.4800 0.2400 0.5400 ;
        RECT 0.0750 0.1875 0.1350 0.2475 ;
        RECT 0.0750 0.8325 0.1350 0.8925 ;
        LAYER M1 ;
        RECT 1.0425 0.4575 1.7400 0.5325 ;
        RECT 1.5225 0.1950 1.6275 0.3825 ;
        RECT 1.5375 0.6225 1.6125 0.8325 ;
        RECT 1.1925 0.6225 1.5375 0.7125 ;
        RECT 1.2075 0.2925 1.5225 0.3825 ;
        RECT 1.1025 0.1950 1.2075 0.3825 ;
        RECT 1.1175 0.6225 1.1925 0.8325 ;
        RECT 0.9675 0.4575 1.0425 0.7875 ;
        RECT 0.3675 0.7125 0.9675 0.7875 ;
        RECT 0.3825 0.1500 0.7725 0.2325 ;
        RECT 0.5400 0.4575 0.7050 0.6375 ;
        RECT 0.3675 0.4575 0.5400 0.5625 ;
        RECT 0.2625 0.7125 0.3675 0.9000 ;
        LAYER VIA1 ;
        RECT 0.9675 0.5025 1.0425 0.5775 ;
        RECT 0.6525 0.1575 0.7275 0.2325 ;
        LAYER M2 ;
        RECT 0.9525 0.2625 1.0575 0.6225 ;
        RECT 0.7725 0.2625 0.9525 0.3375 ;
        RECT 0.6975 0.1575 0.7725 0.3375 ;
        RECT 0.6075 0.1575 0.6975 0.2325 ;
    END
END AN2_0111


MACRO AN2_1000
    CLASS CORE ;
    FOREIGN AN2_1000 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.8400 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.7275 0.1500 0.8025 0.9000 ;
        RECT 0.6975 0.1500 0.7275 0.3825 ;
        RECT 0.6975 0.6675 0.7275 0.9000 ;
        END
    END Z
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.1875 0.2625 0.6525 0.3375 ;
        VIA 0.4800 0.3000 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.4575 0.8625 0.6075 0.9375 ;
        RECT 0.3825 0.4125 0.4575 0.9375 ;
        RECT 0.1875 0.4125 0.3825 0.4875 ;
        RECT 0.0675 0.8625 0.3825 0.9375 ;
        VIA 0.2700 0.4500 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.5925 -0.0750 0.8400 0.0750 ;
        RECT 0.4575 -0.0750 0.5925 0.1800 ;
        RECT 0.0000 -0.0750 0.4575 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.6000 0.9750 0.8400 1.1250 ;
        RECT 0.4650 0.8550 0.6000 1.1250 ;
        RECT 0.1650 0.9750 0.4650 1.1250 ;
        RECT 0.0450 0.8250 0.1650 1.1250 ;
        RECT 0.0000 0.9750 0.0450 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 0.7050 0.1800 0.7650 0.2400 ;
        RECT 0.7050 0.8025 0.7650 0.8625 ;
        RECT 0.5925 0.4950 0.6525 0.5550 ;
        RECT 0.4950 0.1200 0.5550 0.1800 ;
        RECT 0.4950 0.8550 0.5550 0.9150 ;
        RECT 0.3975 0.4800 0.4575 0.5400 ;
        RECT 0.2850 0.8175 0.3450 0.8775 ;
        RECT 0.1875 0.4800 0.2475 0.5400 ;
        RECT 0.0750 0.1575 0.1350 0.2175 ;
        RECT 0.0750 0.8325 0.1350 0.8925 ;
        LAYER M1 ;
        RECT 0.6225 0.4650 0.6525 0.5850 ;
        RECT 0.5475 0.4650 0.6225 0.7500 ;
        RECT 0.4725 0.2550 0.5625 0.3450 ;
        RECT 0.3675 0.6750 0.5475 0.7500 ;
        RECT 0.3975 0.2550 0.4725 0.5700 ;
        RECT 0.2625 0.6750 0.3675 0.9000 ;
        RECT 0.1875 0.3375 0.3225 0.6000 ;
        RECT 0.1125 0.6750 0.2625 0.7500 ;
        RECT 0.1125 0.1500 0.1650 0.2250 ;
        RECT 0.0375 0.1500 0.1125 0.7500 ;
    END
END AN2_1000


MACRO AN2_1010
    CLASS CORE ;
    FOREIGN AN2_1010 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.8400 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.7275 0.2175 0.8025 0.8325 ;
        RECT 0.6975 0.2175 0.7275 0.3825 ;
        RECT 0.6975 0.6675 0.7275 0.8325 ;
        END
    END Z
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.4725 0.2550 0.5625 0.3450 ;
        RECT 0.3975 0.2550 0.4725 0.5700 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.2475 0.2175 0.3225 0.6000 ;
        RECT 0.1875 0.3375 0.2475 0.6000 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.5925 -0.0750 0.8400 0.0750 ;
        RECT 0.4575 -0.0750 0.5925 0.1800 ;
        RECT 0.0000 -0.0750 0.4575 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.6000 0.9750 0.8400 1.1250 ;
        RECT 0.4650 0.8550 0.6000 1.1250 ;
        RECT 0.1650 0.9750 0.4650 1.1250 ;
        RECT 0.0450 0.8250 0.1650 1.1250 ;
        RECT 0.0000 0.9750 0.0450 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 0.7050 0.2625 0.7650 0.3225 ;
        RECT 0.7050 0.7275 0.7650 0.7875 ;
        RECT 0.5925 0.4950 0.6525 0.5550 ;
        RECT 0.4950 0.1200 0.5550 0.1800 ;
        RECT 0.4950 0.8550 0.5550 0.9150 ;
        RECT 0.3975 0.4800 0.4575 0.5400 ;
        RECT 0.2850 0.8175 0.3450 0.8775 ;
        RECT 0.1875 0.4800 0.2475 0.5400 ;
        RECT 0.0750 0.1725 0.1350 0.2325 ;
        RECT 0.0750 0.8325 0.1350 0.8925 ;
        LAYER M1 ;
        RECT 0.6225 0.4650 0.6525 0.5850 ;
        RECT 0.5475 0.4650 0.6225 0.7500 ;
        RECT 0.3675 0.6750 0.5475 0.7500 ;
        RECT 0.2625 0.6750 0.3675 0.9000 ;
        RECT 0.1125 0.6750 0.2625 0.7500 ;
        RECT 0.1125 0.1500 0.1650 0.2550 ;
        RECT 0.0375 0.1500 0.1125 0.7500 ;
    END
END AN2_1010


MACRO AN3_0011
    CLASS CORE ;
    FOREIGN AN3_0011 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.2600 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 1.1475 0.3150 1.2225 0.7350 ;
        RECT 0.9825 0.3150 1.1475 0.3900 ;
        RECT 0.9825 0.6600 1.1475 0.7350 ;
        RECT 0.9075 0.2175 0.9825 0.3900 ;
        RECT 0.9075 0.6600 0.9825 0.8325 ;
        END
    END Z
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.3525 0.5625 0.8175 0.6375 ;
        VIA 0.6000 0.6000 VIA12_square ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.2325 0.4125 0.6975 0.4875 ;
        VIA 0.3975 0.4500 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.1575 0.2625 0.6225 0.3375 ;
        VIA 0.2475 0.3000 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.2150 -0.0750 1.2600 0.0750 ;
        RECT 1.0950 -0.0750 1.2150 0.2400 ;
        RECT 0.7950 -0.0750 1.0950 0.0750 ;
        RECT 0.6750 -0.0750 0.7950 0.2400 ;
        RECT 0.0000 -0.0750 0.6750 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.2150 0.9750 1.2600 1.1250 ;
        RECT 1.0950 0.8100 1.2150 1.1250 ;
        RECT 0.7950 0.9750 1.0950 1.1250 ;
        RECT 0.6750 0.8700 0.7950 1.1250 ;
        RECT 0.3750 0.9750 0.6750 1.1250 ;
        RECT 0.2550 0.8700 0.3750 1.1250 ;
        RECT 0.0000 0.9750 0.2550 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.1250 0.1575 1.1850 0.2175 ;
        RECT 1.1250 0.8325 1.1850 0.8925 ;
        RECT 1.0125 0.4950 1.0725 0.5550 ;
        RECT 0.9150 0.2475 0.9750 0.3075 ;
        RECT 0.9150 0.7125 0.9750 0.7725 ;
        RECT 0.8100 0.4950 0.8700 0.5550 ;
        RECT 0.7050 0.1575 0.7650 0.2175 ;
        RECT 0.7050 0.8700 0.7650 0.9300 ;
        RECT 0.6000 0.4875 0.6600 0.5475 ;
        RECT 0.4950 0.8175 0.5550 0.8775 ;
        RECT 0.3825 0.4875 0.4425 0.5475 ;
        RECT 0.2850 0.8700 0.3450 0.9300 ;
        RECT 0.1875 0.4875 0.2475 0.5475 ;
        RECT 0.0750 0.2100 0.1350 0.2700 ;
        RECT 0.0750 0.8175 0.1350 0.8775 ;
        LAYER M1 ;
        RECT 0.8325 0.4650 1.0725 0.5850 ;
        RECT 0.7575 0.4650 0.8325 0.7950 ;
        RECT 0.5850 0.7200 0.7575 0.7950 ;
        RECT 0.5175 0.4050 0.6825 0.6450 ;
        RECT 0.4650 0.7200 0.5850 0.9000 ;
        RECT 0.1575 0.7200 0.4650 0.7950 ;
        RECT 0.3600 0.2175 0.4425 0.6150 ;
        RECT 0.2100 0.2175 0.2850 0.6150 ;
        RECT 0.1875 0.4275 0.2100 0.6150 ;
        RECT 0.1125 0.7200 0.1575 0.9000 ;
        RECT 0.1125 0.1800 0.1350 0.3000 ;
        RECT 0.0525 0.1800 0.1125 0.9000 ;
        RECT 0.0375 0.1800 0.0525 0.7950 ;
    END
END AN3_0011


MACRO AN3_0100
    CLASS CORE ;
    FOREIGN AN3_0100 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.7800 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 2.9925 0.2775 3.1500 0.3975 ;
        RECT 2.9925 0.6225 3.1500 0.7425 ;
        RECT 2.6775 0.2775 2.9925 0.7425 ;
        RECT 2.5200 0.2775 2.6775 0.3975 ;
        RECT 2.5200 0.6225 2.6775 0.7425 ;
        VIA 2.9925 0.3375 VIA12_slot ;
        VIA 2.9925 0.6825 VIA12_slot ;
        VIA 2.6775 0.3375 VIA12_slot ;
        VIA 2.6775 0.6825 VIA12_slot ;
        END
    END Z
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.5375 0.4125 2.0025 0.4875 ;
        VIA 1.8450 0.4500 VIA12_square ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.1925 0.5625 1.4325 0.6375 ;
        RECT 1.1175 0.4125 1.1925 0.6375 ;
        RECT 0.8625 0.4125 1.1175 0.4875 ;
        VIA 1.1550 0.5100 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.6300 0.5625 0.8700 0.6375 ;
        RECT 0.5550 0.4125 0.6300 0.6375 ;
        RECT 0.3150 0.4125 0.5550 0.4875 ;
        VIA 0.5925 0.5100 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 3.7275 -0.0750 3.7800 0.0750 ;
        RECT 3.6225 -0.0750 3.7275 0.3075 ;
        RECT 3.3150 -0.0750 3.6225 0.0750 ;
        RECT 3.1950 -0.0750 3.3150 0.2025 ;
        RECT 2.8950 -0.0750 3.1950 0.0750 ;
        RECT 2.7750 -0.0750 2.8950 0.2025 ;
        RECT 2.4750 -0.0750 2.7750 0.0750 ;
        RECT 2.3550 -0.0750 2.4750 0.2025 ;
        RECT 2.0325 -0.0750 2.3550 0.0750 ;
        RECT 1.9575 -0.0750 2.0325 0.3075 ;
        RECT 1.6350 -0.0750 1.9575 0.0750 ;
        RECT 1.5150 -0.0750 1.6350 0.1875 ;
        RECT 0.0000 -0.0750 1.5150 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 3.7275 0.9750 3.7800 1.1250 ;
        RECT 3.6225 0.6450 3.7275 1.1250 ;
        RECT 3.3150 0.9750 3.6225 1.1250 ;
        RECT 3.1950 0.8250 3.3150 1.1250 ;
        RECT 2.8950 0.9750 3.1950 1.1250 ;
        RECT 2.7750 0.8250 2.8950 1.1250 ;
        RECT 2.4750 0.9750 2.7750 1.1250 ;
        RECT 2.3550 0.8250 2.4750 1.1250 ;
        RECT 2.0475 0.9750 2.3550 1.1250 ;
        RECT 1.9425 0.8100 2.0475 1.1250 ;
        RECT 1.6275 0.9750 1.9425 1.1250 ;
        RECT 1.5225 0.8100 1.6275 1.1250 ;
        RECT 1.2075 0.9750 1.5225 1.1250 ;
        RECT 1.1025 0.8100 1.2075 1.1250 ;
        RECT 0.7875 0.9750 1.1025 1.1250 ;
        RECT 0.6825 0.8100 0.7875 1.1250 ;
        RECT 0.3675 0.9750 0.6825 1.1250 ;
        RECT 0.2625 0.8100 0.3675 1.1250 ;
        RECT 0.0000 0.9750 0.2625 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 3.6450 0.2175 3.7050 0.2775 ;
        RECT 3.6450 0.6675 3.7050 0.7275 ;
        RECT 3.6450 0.8325 3.7050 0.8925 ;
        RECT 3.5400 0.4800 3.6000 0.5400 ;
        RECT 3.4350 0.3075 3.4950 0.3675 ;
        RECT 3.4350 0.6525 3.4950 0.7125 ;
        RECT 3.3300 0.4800 3.3900 0.5400 ;
        RECT 3.2250 0.1350 3.2850 0.1950 ;
        RECT 3.2250 0.8325 3.2850 0.8925 ;
        RECT 3.1200 0.4800 3.1800 0.5400 ;
        RECT 3.0150 0.3075 3.0750 0.3675 ;
        RECT 3.0150 0.6525 3.0750 0.7125 ;
        RECT 2.9100 0.4800 2.9700 0.5400 ;
        RECT 2.8050 0.1350 2.8650 0.1950 ;
        RECT 2.8050 0.8325 2.8650 0.8925 ;
        RECT 2.7000 0.4800 2.7600 0.5400 ;
        RECT 2.5950 0.3075 2.6550 0.3675 ;
        RECT 2.5950 0.6525 2.6550 0.7125 ;
        RECT 2.4900 0.4800 2.5500 0.5400 ;
        RECT 2.3850 0.1350 2.4450 0.1950 ;
        RECT 2.3850 0.8325 2.4450 0.8925 ;
        RECT 2.2800 0.4800 2.3400 0.5400 ;
        RECT 2.1750 0.3075 2.2350 0.3675 ;
        RECT 2.1750 0.6525 2.2350 0.7125 ;
        RECT 2.0700 0.4800 2.1300 0.5400 ;
        RECT 1.9650 0.2175 2.0250 0.2775 ;
        RECT 1.9650 0.8325 2.0250 0.8925 ;
        RECT 1.8600 0.4800 1.9200 0.5400 ;
        RECT 1.7550 0.2700 1.8150 0.3300 ;
        RECT 1.7550 0.6675 1.8150 0.7275 ;
        RECT 1.6500 0.4800 1.7100 0.5400 ;
        RECT 1.5450 0.1200 1.6050 0.1800 ;
        RECT 1.5450 0.8325 1.6050 0.8925 ;
        RECT 1.4400 0.4800 1.5000 0.5400 ;
        RECT 1.3350 0.3075 1.3950 0.3675 ;
        RECT 1.3350 0.6675 1.3950 0.7275 ;
        RECT 1.2300 0.4800 1.2900 0.5400 ;
        RECT 1.1250 0.1575 1.1850 0.2175 ;
        RECT 1.1250 0.8325 1.1850 0.8925 ;
        RECT 1.0200 0.4800 1.0800 0.5400 ;
        RECT 0.9150 0.3075 0.9750 0.3675 ;
        RECT 0.9150 0.6675 0.9750 0.7275 ;
        RECT 0.8100 0.4800 0.8700 0.5400 ;
        RECT 0.7050 0.1575 0.7650 0.2175 ;
        RECT 0.7050 0.8325 0.7650 0.8925 ;
        RECT 0.6000 0.4800 0.6600 0.5400 ;
        RECT 0.4950 0.3075 0.5550 0.3675 ;
        RECT 0.4950 0.6675 0.5550 0.7275 ;
        RECT 0.3900 0.4800 0.4500 0.5400 ;
        RECT 0.2850 0.1575 0.3450 0.2175 ;
        RECT 0.2850 0.8325 0.3450 0.8925 ;
        RECT 0.1875 0.4800 0.2475 0.5400 ;
        RECT 0.0750 0.3075 0.1350 0.3675 ;
        RECT 0.0750 0.6675 0.1350 0.7275 ;
        LAYER M1 ;
        RECT 2.0775 0.4725 3.6300 0.5475 ;
        RECT 2.1525 0.2775 3.5250 0.3975 ;
        RECT 2.1525 0.6225 3.5250 0.7425 ;
        RECT 2.0025 0.4725 2.0775 0.7350 ;
        RECT 0.1125 0.6600 2.0025 0.7350 ;
        RECT 1.7625 0.4125 1.9275 0.5700 ;
        RECT 1.5225 0.2625 1.8450 0.3375 ;
        RECT 1.4325 0.4500 1.7625 0.5700 ;
        RECT 1.4475 0.2625 1.5225 0.3750 ;
        RECT 0.8850 0.3000 1.4475 0.3750 ;
        RECT 0.8025 0.4500 1.2975 0.5700 ;
        RECT 0.2550 0.1500 1.2150 0.2250 ;
        RECT 0.1875 0.4500 0.6750 0.5700 ;
        RECT 0.1125 0.3000 0.5850 0.3750 ;
        RECT 0.0375 0.3000 0.1125 0.7350 ;
        LAYER M2 ;
        RECT 3.0225 0.2775 3.1500 0.3975 ;
        RECT 3.0225 0.6225 3.1500 0.7425 ;
        RECT 2.5200 0.2775 2.6475 0.3975 ;
        RECT 2.5200 0.6225 2.6475 0.7425 ;
    END
END AN3_0100


MACRO AN3_0111
    CLASS CORE ;
    FOREIGN AN3_0111 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.3100 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 1.6275 0.2550 1.9425 0.7650 ;
        VIA 1.7850 0.3375 VIA12_slot ;
        VIA 1.7850 0.6825 VIA12_slot ;
        END
    END Z
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.1625 0.4125 1.2675 0.5775 ;
        RECT 0.1725 0.4125 1.1625 0.4875 ;
        VIA 1.2150 0.4950 VIA12_square ;
        VIA 0.2550 0.4500 VIA12_square ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.3525 0.2625 0.8175 0.3375 ;
        VIA 0.4950 0.3000 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.4425 0.5625 0.9075 0.6375 ;
        VIA 0.8100 0.6000 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 2.2575 -0.0750 2.3100 0.0750 ;
        RECT 2.1525 -0.0750 2.2575 0.3075 ;
        RECT 1.8450 -0.0750 2.1525 0.0750 ;
        RECT 1.7250 -0.0750 1.8450 0.2025 ;
        RECT 1.4250 -0.0750 1.7250 0.0750 ;
        RECT 1.3050 -0.0750 1.4250 0.1875 ;
        RECT 0.1425 -0.0750 1.3050 0.0750 ;
        RECT 0.0675 -0.0750 0.1425 0.3075 ;
        RECT 0.0000 -0.0750 0.0675 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 2.2575 0.9750 2.3100 1.1250 ;
        RECT 2.1525 0.6450 2.2575 1.1250 ;
        RECT 1.8450 0.9750 2.1525 1.1250 ;
        RECT 1.7250 0.8250 1.8450 1.1250 ;
        RECT 1.4250 0.9750 1.7250 1.1250 ;
        RECT 1.3050 0.8625 1.4250 1.1250 ;
        RECT 1.0050 0.9750 1.3050 1.1250 ;
        RECT 0.8850 0.8625 1.0050 1.1250 ;
        RECT 0.5850 0.9750 0.8850 1.1250 ;
        RECT 0.4650 0.8625 0.5850 1.1250 ;
        RECT 0.1425 0.9750 0.4650 1.1250 ;
        RECT 0.0675 0.6375 0.1425 1.1250 ;
        RECT 0.0000 0.9750 0.0675 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 2.1750 0.2175 2.2350 0.2775 ;
        RECT 2.1750 0.6675 2.2350 0.7275 ;
        RECT 2.1750 0.8325 2.2350 0.8925 ;
        RECT 2.0700 0.4800 2.1300 0.5400 ;
        RECT 1.9650 0.3075 2.0250 0.3675 ;
        RECT 1.9650 0.6525 2.0250 0.7125 ;
        RECT 1.8600 0.4800 1.9200 0.5400 ;
        RECT 1.7550 0.1350 1.8150 0.1950 ;
        RECT 1.7550 0.8325 1.8150 0.8925 ;
        RECT 1.6500 0.4800 1.7100 0.5400 ;
        RECT 1.5450 0.3075 1.6050 0.3675 ;
        RECT 1.5450 0.6525 1.6050 0.7125 ;
        RECT 1.4400 0.4800 1.5000 0.5400 ;
        RECT 1.3350 0.1275 1.3950 0.1875 ;
        RECT 1.3350 0.8700 1.3950 0.9300 ;
        RECT 1.2300 0.4800 1.2900 0.5400 ;
        RECT 1.1250 0.7200 1.1850 0.7800 ;
        RECT 0.7050 0.7200 0.7650 0.7800 ;
        RECT 0.6000 0.4950 0.6600 0.5550 ;
        RECT 0.4950 0.8700 0.5550 0.9300 ;
        RECT 0.3900 0.4875 0.4500 0.5475 ;
        RECT 0.2850 0.7200 0.3450 0.7800 ;
        RECT 0.1800 0.4650 0.2400 0.5250 ;
        RECT 0.0750 0.2175 0.1350 0.2775 ;
        RECT 0.0750 0.6675 0.1350 0.7275 ;
        RECT 0.0750 0.8325 0.1350 0.8925 ;
        RECT 1.0200 0.4875 1.0800 0.5475 ;
        RECT 0.9150 0.8700 0.9750 0.9300 ;
        RECT 0.8100 0.4950 0.8700 0.5550 ;
        RECT 0.7050 0.1650 0.7650 0.2250 ;
        LAYER M1 ;
        RECT 1.4475 0.4725 2.1600 0.5475 ;
        RECT 1.5225 0.2775 2.0550 0.3975 ;
        RECT 1.5225 0.6225 2.0550 0.7425 ;
        RECT 1.3725 0.2625 1.4475 0.7875 ;
        RECT 1.2225 0.2625 1.3725 0.3375 ;
        RECT 0.2550 0.7125 1.3725 0.7875 ;
        RECT 1.1550 0.4125 1.2975 0.6375 ;
        RECT 1.1475 0.1575 1.2225 0.3375 ;
        RECT 0.6750 0.1575 1.1475 0.2325 ;
        RECT 1.0425 0.4500 1.0800 0.5850 ;
        RECT 0.9675 0.3225 1.0425 0.5850 ;
        RECT 0.5625 0.3225 0.9675 0.3975 ;
        RECT 0.7275 0.4725 0.8925 0.6375 ;
        RECT 0.5775 0.4725 0.7275 0.5775 ;
        RECT 0.5025 0.2175 0.5625 0.3975 ;
        RECT 0.4275 0.2175 0.5025 0.5700 ;
        RECT 0.3675 0.4650 0.4275 0.5700 ;
        RECT 0.2175 0.2250 0.2925 0.5325 ;
        RECT 0.1350 0.4350 0.2175 0.5325 ;
    END
END AN3_0111


MACRO AN3_1000
    CLASS CORE ;
    FOREIGN AN3_1000 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.0500 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.9375 0.1500 1.0125 0.9000 ;
        RECT 0.9075 0.1500 0.9375 0.3150 ;
        RECT 0.9075 0.6675 0.9375 0.9000 ;
        END
    END Z
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.3525 0.5625 0.8175 0.6375 ;
        VIA 0.6000 0.6000 VIA12_square ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.2325 0.4125 0.6975 0.4875 ;
        VIA 0.4050 0.4500 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.1575 0.2625 0.6225 0.3375 ;
        VIA 0.2550 0.3000 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.7950 -0.0750 1.0500 0.0750 ;
        RECT 0.6750 -0.0750 0.7950 0.1800 ;
        RECT 0.0000 -0.0750 0.6750 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.7950 0.9750 1.0500 1.1250 ;
        RECT 0.6750 0.8700 0.7950 1.1250 ;
        RECT 0.3750 0.9750 0.6750 1.1250 ;
        RECT 0.2550 0.8700 0.3750 1.1250 ;
        RECT 0.0000 0.9750 0.2550 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 0.9150 0.1800 0.9750 0.2400 ;
        RECT 0.9150 0.8100 0.9750 0.8700 ;
        RECT 0.8025 0.4875 0.8625 0.5475 ;
        RECT 0.7050 0.1200 0.7650 0.1800 ;
        RECT 0.7050 0.8700 0.7650 0.9300 ;
        RECT 0.6000 0.4875 0.6600 0.5475 ;
        RECT 0.4950 0.8175 0.5550 0.8775 ;
        RECT 0.3825 0.5250 0.4425 0.5850 ;
        RECT 0.2850 0.8700 0.3450 0.9300 ;
        RECT 0.1875 0.5100 0.2475 0.5700 ;
        RECT 0.0750 0.1800 0.1350 0.2400 ;
        RECT 0.0750 0.8175 0.1350 0.8775 ;
        LAYER M1 ;
        RECT 0.8325 0.4575 0.8625 0.5775 ;
        RECT 0.7575 0.4575 0.8325 0.7950 ;
        RECT 0.5850 0.7200 0.7575 0.7950 ;
        RECT 0.5250 0.4050 0.6825 0.6450 ;
        RECT 0.4650 0.7200 0.5850 0.9000 ;
        RECT 0.5175 0.5400 0.5250 0.6450 ;
        RECT 0.1575 0.7200 0.4650 0.7950 ;
        RECT 0.4425 0.2175 0.4500 0.4875 ;
        RECT 0.3675 0.2175 0.4425 0.6150 ;
        RECT 0.2175 0.2175 0.2925 0.6150 ;
        RECT 0.1875 0.4275 0.2175 0.6150 ;
        RECT 0.1125 0.7200 0.1575 0.9000 ;
        RECT 0.1125 0.1500 0.1425 0.2700 ;
        RECT 0.0525 0.1500 0.1125 0.9000 ;
        RECT 0.0375 0.1500 0.0525 0.7950 ;
    END
END AN3_1000


MACRO AN3_1010
    CLASS CORE ;
    FOREIGN AN3_1010 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.0500 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.9375 0.2175 1.0125 0.8325 ;
        RECT 0.9075 0.2175 0.9375 0.3825 ;
        RECT 0.9075 0.6675 0.9375 0.8325 ;
        END
    END Z
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.5175 0.4050 0.6825 0.6450 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.3600 0.2175 0.4425 0.6150 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.2100 0.2175 0.2850 0.6150 ;
        RECT 0.1875 0.4275 0.2100 0.6150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.7950 -0.0750 1.0500 0.0750 ;
        RECT 0.6750 -0.0750 0.7950 0.2850 ;
        RECT 0.0000 -0.0750 0.6750 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.7950 0.9750 1.0500 1.1250 ;
        RECT 0.6750 0.8700 0.7950 1.1250 ;
        RECT 0.3750 0.9750 0.6750 1.1250 ;
        RECT 0.2550 0.8700 0.3750 1.1250 ;
        RECT 0.0000 0.9750 0.2550 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 0.9150 0.2475 0.9750 0.3075 ;
        RECT 0.9150 0.7125 0.9750 0.7725 ;
        RECT 0.8025 0.4875 0.8625 0.5475 ;
        RECT 0.7050 0.2100 0.7650 0.2700 ;
        RECT 0.7050 0.8700 0.7650 0.9300 ;
        RECT 0.6000 0.4875 0.6600 0.5475 ;
        RECT 0.4950 0.8175 0.5550 0.8775 ;
        RECT 0.3825 0.5250 0.4425 0.5850 ;
        RECT 0.2850 0.8700 0.3450 0.9300 ;
        RECT 0.1875 0.5100 0.2475 0.5700 ;
        RECT 0.0750 0.2100 0.1350 0.2700 ;
        RECT 0.0750 0.8175 0.1350 0.8775 ;
        LAYER M1 ;
        RECT 0.8325 0.4575 0.8625 0.5775 ;
        RECT 0.7575 0.4575 0.8325 0.7950 ;
        RECT 0.5850 0.7200 0.7575 0.7950 ;
        RECT 0.4650 0.7200 0.5850 0.9000 ;
        RECT 0.1575 0.7200 0.4650 0.7950 ;
        RECT 0.1125 0.7200 0.1575 0.9000 ;
        RECT 0.1125 0.1800 0.1350 0.3000 ;
        RECT 0.0525 0.1800 0.1125 0.9000 ;
        RECT 0.0375 0.1800 0.0525 0.7950 ;
    END
END AN3_1010


MACRO AN4_0011
    CLASS CORE ;
    FOREIGN AN4_0011 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.4700 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 1.3575 0.3075 1.4325 0.7425 ;
        RECT 1.1925 0.3075 1.3575 0.3825 ;
        RECT 1.1925 0.6675 1.3575 0.7425 ;
        RECT 1.1175 0.2175 1.1925 0.3825 ;
        RECT 1.1175 0.6675 1.1925 0.8550 ;
        END
    END Z
    PIN A4
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.7275 0.4125 1.1925 0.4875 ;
        VIA 0.8100 0.4500 VIA12_square ;
        END
    END A4
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.5550 0.2625 0.6900 0.3375 ;
        RECT 0.4800 0.2625 0.5550 0.4275 ;
        RECT 0.1500 0.2625 0.4800 0.3375 ;
        VIA 0.5175 0.3450 VIA12_square ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.4275 0.7125 0.8925 0.7875 ;
        RECT 0.3525 0.5250 0.4275 0.7875 ;
        VIA 0.3900 0.6075 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1425 0.4650 0.2325 0.5850 ;
        RECT 0.0675 0.3675 0.1425 0.6825 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.4250 -0.0750 1.4700 0.0750 ;
        RECT 1.3050 -0.0750 1.4250 0.2175 ;
        RECT 1.0050 -0.0750 1.3050 0.0750 ;
        RECT 0.8850 -0.0750 1.0050 0.1800 ;
        RECT 0.0000 -0.0750 0.8850 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.4250 0.9750 1.4700 1.1250 ;
        RECT 1.3050 0.8175 1.4250 1.1250 ;
        RECT 1.0050 0.9750 1.3050 1.1250 ;
        RECT 0.8850 0.8700 1.0050 1.1250 ;
        RECT 0.5850 0.9750 0.8850 1.1250 ;
        RECT 0.4650 0.8700 0.5850 1.1250 ;
        RECT 0.1650 0.9750 0.4650 1.1250 ;
        RECT 0.0450 0.8250 0.1650 1.1250 ;
        RECT 0.0000 0.9750 0.0450 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.3350 0.1575 1.3950 0.2175 ;
        RECT 1.3350 0.8325 1.3950 0.8925 ;
        RECT 1.2225 0.4950 1.2825 0.5550 ;
        RECT 1.1250 0.2475 1.1850 0.3075 ;
        RECT 1.1250 0.7650 1.1850 0.8250 ;
        RECT 1.0200 0.4950 1.0800 0.5550 ;
        RECT 0.9150 0.1200 0.9750 0.1800 ;
        RECT 0.9150 0.8700 0.9750 0.9300 ;
        RECT 0.8100 0.4650 0.8700 0.5250 ;
        RECT 0.7050 0.8250 0.7650 0.8850 ;
        RECT 0.5925 0.4875 0.6525 0.5475 ;
        RECT 0.4950 0.8700 0.5550 0.9300 ;
        RECT 0.3900 0.4950 0.4500 0.5550 ;
        RECT 0.2850 0.7950 0.3450 0.8550 ;
        RECT 0.1725 0.4950 0.2325 0.5550 ;
        RECT 0.0750 0.1650 0.1350 0.2250 ;
        RECT 0.0750 0.8325 0.1350 0.8925 ;
        LAYER M1 ;
        RECT 1.0425 0.4650 1.2825 0.5850 ;
        RECT 0.9675 0.2625 1.0425 0.7950 ;
        RECT 0.8100 0.2625 0.9675 0.3375 ;
        RECT 0.7950 0.7200 0.9675 0.7950 ;
        RECT 0.7275 0.4125 0.8925 0.6450 ;
        RECT 0.7350 0.1500 0.8100 0.3375 ;
        RECT 0.6750 0.7200 0.7950 0.9000 ;
        RECT 0.1500 0.1500 0.7350 0.2250 ;
        RECT 0.3675 0.7200 0.6750 0.7950 ;
        RECT 0.5775 0.3075 0.6525 0.6150 ;
        RECT 0.4275 0.3075 0.5775 0.3825 ;
        RECT 0.3075 0.4575 0.5025 0.6450 ;
        RECT 0.2400 0.7200 0.3675 0.8850 ;
        RECT 0.0450 0.1500 0.1500 0.2550 ;
    END
END AN4_0011


MACRO AN4_0100
    CLASS CORE ;
    FOREIGN AN4_0100 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.4100 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 3.6225 0.2775 3.7800 0.3975 ;
        RECT 3.6225 0.6225 3.7800 0.7425 ;
        RECT 3.3075 0.2775 3.6225 0.7425 ;
        RECT 3.1500 0.2775 3.3075 0.3975 ;
        RECT 3.1500 0.6225 3.3075 0.7425 ;
        VIA 3.6225 0.3375 VIA12_slot ;
        VIA 3.6225 0.6825 VIA12_slot ;
        VIA 3.3075 0.3375 VIA12_slot ;
        VIA 3.3075 0.6825 VIA12_slot ;
        END
    END Z
    PIN A4
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 2.4525 0.5625 2.6925 0.6375 ;
        RECT 2.3775 0.4125 2.4525 0.6375 ;
        RECT 2.1375 0.4125 2.3775 0.4875 ;
        VIA 2.4150 0.5025 VIA12_square ;
        END
    END A4
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.8225 0.5625 2.0625 0.6375 ;
        RECT 1.7475 0.4125 1.8225 0.6375 ;
        RECT 1.5075 0.4125 1.7475 0.4875 ;
        VIA 1.7850 0.5100 VIA12_square ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.1925 0.5625 1.4325 0.6375 ;
        RECT 1.1175 0.4125 1.1925 0.6375 ;
        RECT 0.8775 0.4125 1.1175 0.4875 ;
        VIA 1.1550 0.5100 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.6375 0.5625 0.8775 0.6375 ;
        RECT 0.5625 0.4125 0.6375 0.6375 ;
        RECT 0.3225 0.4125 0.5625 0.4875 ;
        VIA 0.6000 0.5100 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 4.3575 -0.0750 4.4100 0.0750 ;
        RECT 4.2525 -0.0750 4.3575 0.3075 ;
        RECT 3.9450 -0.0750 4.2525 0.0750 ;
        RECT 3.8250 -0.0750 3.9450 0.2025 ;
        RECT 3.5250 -0.0750 3.8250 0.0750 ;
        RECT 3.4050 -0.0750 3.5250 0.2025 ;
        RECT 3.1050 -0.0750 3.4050 0.0750 ;
        RECT 2.9850 -0.0750 3.1050 0.2025 ;
        RECT 2.6625 -0.0750 2.9850 0.0750 ;
        RECT 2.5875 -0.0750 2.6625 0.3075 ;
        RECT 2.2575 -0.0750 2.5875 0.0750 ;
        RECT 2.1525 -0.0750 2.2575 0.2250 ;
        RECT 0.0000 -0.0750 2.1525 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 4.3575 0.9750 4.4100 1.1250 ;
        RECT 4.2525 0.6450 4.3575 1.1250 ;
        RECT 3.9450 0.9750 4.2525 1.1250 ;
        RECT 3.8250 0.8250 3.9450 1.1250 ;
        RECT 3.5250 0.9750 3.8250 1.1250 ;
        RECT 3.4050 0.8250 3.5250 1.1250 ;
        RECT 3.1050 0.9750 3.4050 1.1250 ;
        RECT 2.9850 0.8250 3.1050 1.1250 ;
        RECT 2.6775 0.9750 2.9850 1.1250 ;
        RECT 2.5725 0.8100 2.6775 1.1250 ;
        RECT 2.2575 0.9750 2.5725 1.1250 ;
        RECT 2.1525 0.8100 2.2575 1.1250 ;
        RECT 1.8375 0.9750 2.1525 1.1250 ;
        RECT 1.7325 0.8100 1.8375 1.1250 ;
        RECT 1.4175 0.9750 1.7325 1.1250 ;
        RECT 1.3125 0.8100 1.4175 1.1250 ;
        RECT 0.9975 0.9750 1.3125 1.1250 ;
        RECT 0.8925 0.8100 0.9975 1.1250 ;
        RECT 0.5775 0.9750 0.8925 1.1250 ;
        RECT 0.4725 0.8100 0.5775 1.1250 ;
        RECT 0.1575 0.9750 0.4725 1.1250 ;
        RECT 0.0525 0.8100 0.1575 1.1250 ;
        RECT 0.0000 0.9750 0.0525 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 4.2750 0.2175 4.3350 0.2775 ;
        RECT 4.2750 0.6675 4.3350 0.7275 ;
        RECT 4.2750 0.8325 4.3350 0.8925 ;
        RECT 4.1700 0.4800 4.2300 0.5400 ;
        RECT 4.0650 0.3075 4.1250 0.3675 ;
        RECT 4.0650 0.6525 4.1250 0.7125 ;
        RECT 3.9600 0.4800 4.0200 0.5400 ;
        RECT 3.8550 0.1350 3.9150 0.1950 ;
        RECT 3.8550 0.8325 3.9150 0.8925 ;
        RECT 3.7500 0.4800 3.8100 0.5400 ;
        RECT 3.6450 0.3075 3.7050 0.3675 ;
        RECT 3.6450 0.6525 3.7050 0.7125 ;
        RECT 3.5400 0.4800 3.6000 0.5400 ;
        RECT 3.4350 0.1350 3.4950 0.1950 ;
        RECT 3.4350 0.8325 3.4950 0.8925 ;
        RECT 3.3300 0.4800 3.3900 0.5400 ;
        RECT 3.2250 0.3075 3.2850 0.3675 ;
        RECT 3.2250 0.6525 3.2850 0.7125 ;
        RECT 3.1200 0.4800 3.1800 0.5400 ;
        RECT 3.0150 0.1350 3.0750 0.1950 ;
        RECT 3.0150 0.8325 3.0750 0.8925 ;
        RECT 2.9100 0.4800 2.9700 0.5400 ;
        RECT 2.8050 0.3075 2.8650 0.3675 ;
        RECT 2.8050 0.6525 2.8650 0.7125 ;
        RECT 2.7000 0.4800 2.7600 0.5400 ;
        RECT 2.5950 0.2175 2.6550 0.2775 ;
        RECT 2.5950 0.8325 2.6550 0.8925 ;
        RECT 2.4900 0.4800 2.5500 0.5400 ;
        RECT 2.3850 0.3075 2.4450 0.3675 ;
        RECT 2.3850 0.6675 2.4450 0.7275 ;
        RECT 2.2800 0.4800 2.3400 0.5400 ;
        RECT 2.1750 0.1425 2.2350 0.2025 ;
        RECT 2.1750 0.8325 2.2350 0.8925 ;
        RECT 2.0700 0.4800 2.1300 0.5400 ;
        RECT 1.9650 0.3075 2.0250 0.3675 ;
        RECT 1.9650 0.6675 2.0250 0.7275 ;
        RECT 1.8600 0.4800 1.9200 0.5400 ;
        RECT 1.7550 0.1575 1.8150 0.2175 ;
        RECT 1.7550 0.8325 1.8150 0.8925 ;
        RECT 1.6500 0.4800 1.7100 0.5400 ;
        RECT 1.5450 0.3075 1.6050 0.3675 ;
        RECT 1.5450 0.6675 1.6050 0.7275 ;
        RECT 1.4400 0.4800 1.5000 0.5400 ;
        RECT 1.3350 0.1575 1.3950 0.2175 ;
        RECT 1.3350 0.8325 1.3950 0.8925 ;
        RECT 1.2300 0.4800 1.2900 0.5400 ;
        RECT 1.1250 0.3075 1.1850 0.3675 ;
        RECT 1.1250 0.6675 1.1850 0.7275 ;
        RECT 1.0200 0.4800 1.0800 0.5400 ;
        RECT 0.9150 0.1575 0.9750 0.2175 ;
        RECT 0.9150 0.8325 0.9750 0.8925 ;
        RECT 0.8100 0.4800 0.8700 0.5400 ;
        RECT 0.7050 0.2850 0.7650 0.3450 ;
        RECT 0.7050 0.6675 0.7650 0.7275 ;
        RECT 0.6000 0.4800 0.6600 0.5400 ;
        RECT 0.4950 0.3075 0.5550 0.3675 ;
        RECT 0.4950 0.8325 0.5550 0.8925 ;
        RECT 0.3900 0.4800 0.4500 0.5400 ;
        RECT 0.2850 0.1575 0.3450 0.2175 ;
        RECT 0.2850 0.6675 0.3450 0.7275 ;
        RECT 0.1875 0.4800 0.2475 0.5400 ;
        RECT 0.0750 0.3075 0.1350 0.3675 ;
        RECT 0.0750 0.8325 0.1350 0.8925 ;
        LAYER M1 ;
        RECT 2.7075 0.4725 4.2600 0.5475 ;
        RECT 2.7825 0.6225 4.1550 0.7425 ;
        RECT 2.7825 0.2775 4.1475 0.3975 ;
        RECT 2.6325 0.4725 2.7075 0.7350 ;
        RECT 0.1125 0.6600 2.6325 0.7350 ;
        RECT 2.0625 0.4500 2.5575 0.5700 ;
        RECT 1.5150 0.3000 2.4750 0.3750 ;
        RECT 1.4175 0.4575 1.9425 0.5625 ;
        RECT 0.8850 0.1500 1.8450 0.2250 ;
        RECT 0.7875 0.4575 1.3125 0.5625 ;
        RECT 0.7800 0.3000 1.2150 0.3750 ;
        RECT 0.7050 0.1500 0.7800 0.3750 ;
        RECT 0.2550 0.1500 0.7050 0.2250 ;
        RECT 0.1875 0.4500 0.6825 0.5700 ;
        RECT 0.1125 0.3000 0.6000 0.3750 ;
        RECT 0.0375 0.3000 0.1125 0.7350 ;
        LAYER M2 ;
        RECT 3.6525 0.2775 3.7800 0.3975 ;
        RECT 3.6525 0.6225 3.7800 0.7425 ;
        RECT 3.1500 0.2775 3.2775 0.3975 ;
        RECT 3.1500 0.6225 3.2775 0.7425 ;
    END
END AN4_0100


MACRO AN4_0111
    CLASS CORE ;
    FOREIGN AN4_0111 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.7300 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 2.0475 0.2550 2.3625 0.7650 ;
        VIA 2.2050 0.3375 VIA12_slot ;
        VIA 2.2050 0.6825 VIA12_slot ;
        END
    END Z
    PIN A4
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.6125 0.2700 1.6875 0.5850 ;
        RECT 1.3125 0.2700 1.6125 0.3450 ;
        RECT 1.2375 0.2700 1.3125 0.4875 ;
        RECT 0.1725 0.4125 1.2375 0.4875 ;
        VIA 1.6500 0.4950 VIA12_square ;
        VIA 0.2550 0.4500 VIA12_square ;
        END
    END A4
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.4100 0.4725 1.4850 0.7875 ;
        RECT 0.5325 0.7125 1.4100 0.7875 ;
        RECT 0.4575 0.5625 0.5325 0.7875 ;
        RECT 0.3675 0.5625 0.4575 0.6375 ;
        VIA 1.4475 0.5550 VIA12_square ;
        VIA 0.4500 0.6000 VIA12_square ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.5925 0.2625 1.0575 0.3375 ;
        VIA 0.6750 0.3000 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.7500 0.5625 1.2150 0.6375 ;
        VIA 1.0050 0.6000 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 2.6775 -0.0750 2.7300 0.0750 ;
        RECT 2.5725 -0.0750 2.6775 0.3075 ;
        RECT 2.2650 -0.0750 2.5725 0.0750 ;
        RECT 2.1450 -0.0750 2.2650 0.1950 ;
        RECT 1.8450 -0.0750 2.1450 0.0750 ;
        RECT 1.7250 -0.0750 1.8450 0.1875 ;
        RECT 0.1425 -0.0750 1.7250 0.0750 ;
        RECT 0.0675 -0.0750 0.1425 0.2850 ;
        RECT 0.0000 -0.0750 0.0675 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 2.6775 0.9750 2.7300 1.1250 ;
        RECT 2.5725 0.6450 2.6775 1.1250 ;
        RECT 2.2650 0.9750 2.5725 1.1250 ;
        RECT 2.1450 0.8250 2.2650 1.1250 ;
        RECT 1.8450 0.9750 2.1450 1.1250 ;
        RECT 1.7250 0.8625 1.8450 1.1250 ;
        RECT 1.4250 0.9750 1.7250 1.1250 ;
        RECT 1.3050 0.8625 1.4250 1.1250 ;
        RECT 1.0050 0.9750 1.3050 1.1250 ;
        RECT 0.8850 0.8625 1.0050 1.1250 ;
        RECT 0.5850 0.9750 0.8850 1.1250 ;
        RECT 0.4650 0.8625 0.5850 1.1250 ;
        RECT 0.1425 0.9750 0.4650 1.1250 ;
        RECT 0.0675 0.6375 0.1425 1.1250 ;
        RECT 0.0000 0.9750 0.0675 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 2.5950 0.2175 2.6550 0.2775 ;
        RECT 2.5950 0.6675 2.6550 0.7275 ;
        RECT 2.5950 0.8325 2.6550 0.8925 ;
        RECT 2.4900 0.4800 2.5500 0.5400 ;
        RECT 2.3850 0.3075 2.4450 0.3675 ;
        RECT 2.3850 0.6525 2.4450 0.7125 ;
        RECT 2.2800 0.4800 2.3400 0.5400 ;
        RECT 2.1750 0.1275 2.2350 0.1875 ;
        RECT 2.1750 0.8325 2.2350 0.8925 ;
        RECT 2.0700 0.4800 2.1300 0.5400 ;
        RECT 1.9650 0.3075 2.0250 0.3675 ;
        RECT 1.9650 0.6525 2.0250 0.7125 ;
        RECT 1.8600 0.4800 1.9200 0.5400 ;
        RECT 1.7550 0.1200 1.8150 0.1800 ;
        RECT 1.7550 0.8700 1.8150 0.9300 ;
        RECT 1.6500 0.4800 1.7100 0.5400 ;
        RECT 1.5450 0.7200 1.6050 0.7800 ;
        RECT 1.4400 0.4800 1.5000 0.5400 ;
        RECT 1.3350 0.8700 1.3950 0.9300 ;
        RECT 1.2300 0.4800 1.2900 0.5400 ;
        RECT 1.1250 0.7200 1.1850 0.7800 ;
        RECT 1.0200 0.4875 1.0800 0.5475 ;
        RECT 0.9150 0.1575 0.9750 0.2175 ;
        RECT 0.9150 0.8700 0.9750 0.9300 ;
        RECT 0.8100 0.4875 0.8700 0.5475 ;
        RECT 0.7050 0.7200 0.7650 0.7800 ;
        RECT 0.6075 0.4875 0.6675 0.5475 ;
        RECT 0.4950 0.8700 0.5550 0.9300 ;
        RECT 0.3900 0.4875 0.4500 0.5475 ;
        RECT 0.2850 0.7200 0.3450 0.7800 ;
        RECT 0.1800 0.4650 0.2400 0.5250 ;
        RECT 0.0750 0.6675 0.1350 0.7275 ;
        RECT 0.0750 0.8325 0.1350 0.8925 ;
        RECT 0.0750 0.1950 0.1350 0.2550 ;
        LAYER M1 ;
        RECT 1.8675 0.4725 2.5800 0.5475 ;
        RECT 1.9425 0.2775 2.4750 0.3975 ;
        RECT 1.9425 0.6225 2.4750 0.7425 ;
        RECT 1.7925 0.2625 1.8675 0.7875 ;
        RECT 1.6425 0.2625 1.7925 0.3375 ;
        RECT 0.2550 0.7125 1.7925 0.7875 ;
        RECT 1.5750 0.4125 1.7175 0.6375 ;
        RECT 1.5675 0.1500 1.6425 0.3375 ;
        RECT 0.8850 0.1500 1.5675 0.2250 ;
        RECT 1.4700 0.4125 1.5000 0.6375 ;
        RECT 1.3725 0.3300 1.4700 0.6375 ;
        RECT 1.2375 0.4500 1.2975 0.5700 ;
        RECT 1.1625 0.3075 1.2375 0.5700 ;
        RECT 0.7125 0.3075 1.1625 0.3825 ;
        RECT 0.9225 0.4575 1.0875 0.6375 ;
        RECT 0.8025 0.4575 0.9225 0.5850 ;
        RECT 0.6075 0.2175 0.7125 0.5775 ;
        RECT 0.3675 0.3675 0.5325 0.6375 ;
        RECT 0.2175 0.2550 0.2925 0.6075 ;
        RECT 0.1350 0.4350 0.2175 0.5325 ;
    END
END AN4_0111


MACRO AN4_1000
    CLASS CORE ;
    FOREIGN AN4_1000 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.2600 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 1.1475 0.1500 1.2225 0.9000 ;
        RECT 1.1175 0.1500 1.1475 0.3825 ;
        RECT 1.1175 0.6675 1.1475 0.9000 ;
        END
    END Z
    PIN A4
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.7275 0.4125 1.1925 0.4875 ;
        VIA 0.8100 0.4500 VIA12_square ;
        END
    END A4
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.5550 0.2625 0.9000 0.3375 ;
        RECT 0.4800 0.2625 0.5550 0.4275 ;
        RECT 0.3600 0.2625 0.4800 0.3375 ;
        VIA 0.5175 0.3450 VIA12_square ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.4275 0.7125 0.8925 0.7875 ;
        RECT 0.3525 0.5250 0.4275 0.7875 ;
        VIA 0.3900 0.6075 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1425 0.4650 0.2325 0.5850 ;
        RECT 0.0675 0.3675 0.1425 0.6825 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.0050 -0.0750 1.2600 0.0750 ;
        RECT 0.8850 -0.0750 1.0050 0.1800 ;
        RECT 0.0000 -0.0750 0.8850 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.0050 0.9750 1.2600 1.1250 ;
        RECT 0.8850 0.8700 1.0050 1.1250 ;
        RECT 0.5850 0.9750 0.8850 1.1250 ;
        RECT 0.4650 0.8700 0.5850 1.1250 ;
        RECT 0.1650 0.9750 0.4650 1.1250 ;
        RECT 0.0450 0.8250 0.1650 1.1250 ;
        RECT 0.0000 0.9750 0.0450 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.1250 0.1800 1.1850 0.2400 ;
        RECT 1.1250 0.8100 1.1850 0.8700 ;
        RECT 1.0125 0.4875 1.0725 0.5475 ;
        RECT 0.9150 0.1200 0.9750 0.1800 ;
        RECT 0.9150 0.8700 0.9750 0.9300 ;
        RECT 0.8100 0.4650 0.8700 0.5250 ;
        RECT 0.7050 0.8250 0.7650 0.8850 ;
        RECT 0.5925 0.4875 0.6525 0.5475 ;
        RECT 0.4950 0.8700 0.5550 0.9300 ;
        RECT 0.3900 0.4950 0.4500 0.5550 ;
        RECT 0.2850 0.7950 0.3450 0.8550 ;
        RECT 0.1725 0.4950 0.2325 0.5550 ;
        RECT 0.0750 0.1650 0.1350 0.2250 ;
        RECT 0.0750 0.8325 0.1350 0.8925 ;
        LAYER M1 ;
        RECT 1.0425 0.4575 1.0725 0.5775 ;
        RECT 0.9675 0.2625 1.0425 0.7950 ;
        RECT 0.8100 0.2625 0.9675 0.3375 ;
        RECT 0.7950 0.7200 0.9675 0.7950 ;
        RECT 0.7275 0.4125 0.8925 0.6450 ;
        RECT 0.7350 0.1500 0.8100 0.3375 ;
        RECT 0.6750 0.7200 0.7950 0.9000 ;
        RECT 0.1500 0.1500 0.7350 0.2250 ;
        RECT 0.3675 0.7200 0.6750 0.7950 ;
        RECT 0.5775 0.3075 0.6525 0.6150 ;
        RECT 0.4275 0.3075 0.5775 0.3825 ;
        RECT 0.3075 0.4575 0.5025 0.6450 ;
        RECT 0.2400 0.7200 0.3675 0.8850 ;
        RECT 0.0450 0.1500 0.1500 0.2550 ;
    END
END AN4_1000


MACRO AN4_1010
    CLASS CORE ;
    FOREIGN AN4_1010 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.2600 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 1.1475 0.2175 1.2225 0.8325 ;
        RECT 1.1175 0.2175 1.1475 0.3825 ;
        RECT 1.1175 0.6675 1.1475 0.8325 ;
        END
    END Z
    PIN A4
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.7275 0.4125 0.8925 0.6375 ;
        END
    END A4
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.5700 0.1800 0.6525 0.5775 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.3825 0.1800 0.4725 0.5775 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.2175 0.1800 0.2925 0.5850 ;
        RECT 0.1875 0.4650 0.2175 0.5850 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.0050 -0.0750 1.2600 0.0750 ;
        RECT 0.8850 -0.0750 1.0050 0.1800 ;
        RECT 0.0000 -0.0750 0.8850 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.0050 0.9750 1.2600 1.1250 ;
        RECT 0.8850 0.8700 1.0050 1.1250 ;
        RECT 0.5850 0.9750 0.8850 1.1250 ;
        RECT 0.4650 0.8700 0.5850 1.1250 ;
        RECT 0.1650 0.9750 0.4650 1.1250 ;
        RECT 0.0450 0.8325 0.1650 1.1250 ;
        RECT 0.0000 0.9750 0.0450 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.1250 0.2700 1.1850 0.3300 ;
        RECT 1.1250 0.7275 1.1850 0.7875 ;
        RECT 1.0125 0.4875 1.0725 0.5475 ;
        RECT 0.9150 0.1200 0.9750 0.1800 ;
        RECT 0.9150 0.8700 0.9750 0.9300 ;
        RECT 0.8100 0.4650 0.8700 0.5250 ;
        RECT 0.7050 0.8250 0.7650 0.8850 ;
        RECT 0.5925 0.4875 0.6525 0.5475 ;
        RECT 0.4950 0.8700 0.5550 0.9300 ;
        RECT 0.3900 0.4875 0.4500 0.5475 ;
        RECT 0.2850 0.8175 0.3450 0.8775 ;
        RECT 0.1875 0.4950 0.2475 0.5550 ;
        RECT 0.0750 0.2325 0.1350 0.2925 ;
        RECT 0.0750 0.8325 0.1350 0.8925 ;
        LAYER M1 ;
        RECT 1.0425 0.4575 1.0725 0.5775 ;
        RECT 0.9675 0.4575 1.0425 0.7950 ;
        RECT 0.7950 0.7200 0.9675 0.7950 ;
        RECT 0.6750 0.7200 0.7950 0.9000 ;
        RECT 0.3675 0.7200 0.6750 0.7950 ;
        RECT 0.3300 0.7200 0.3675 0.9000 ;
        RECT 0.2625 0.6825 0.3300 0.9000 ;
        RECT 0.1125 0.6825 0.2625 0.7575 ;
        RECT 0.1125 0.2025 0.1425 0.3225 ;
        RECT 0.0375 0.2025 0.1125 0.7575 ;
    END
END AN4_1010


MACRO AO211_0011
    CLASS CORE ;
    FOREIGN AO211_0011 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.4700 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 1.3575 0.3075 1.4325 0.7425 ;
        RECT 1.1925 0.3075 1.3575 0.3825 ;
        RECT 1.1925 0.6675 1.3575 0.7425 ;
        RECT 1.1175 0.2175 1.1925 0.3825 ;
        RECT 1.1175 0.6675 1.1925 0.8550 ;
        END
    END Z
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.8325 0.6675 0.9075 0.9375 ;
        RECT 0.3675 0.8625 0.8325 0.9375 ;
        VIA 0.8700 0.7500 VIA12_square ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.7275 0.4125 1.1925 0.4875 ;
        RECT 0.6525 0.4125 0.7275 0.6450 ;
        VIA 0.6900 0.5175 VIA12_square ;
        END
    END B
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.4275 0.1125 0.8925 0.1875 ;
        RECT 0.3525 0.1125 0.4275 0.5250 ;
        VIA 0.3900 0.4425 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1725 0.4275 0.2325 0.5700 ;
        RECT 0.1425 0.3525 0.1725 0.5700 ;
        RECT 0.0675 0.3525 0.1425 0.6825 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.4250 -0.0750 1.4700 0.0750 ;
        RECT 1.3050 -0.0750 1.4250 0.2175 ;
        RECT 1.0050 -0.0750 1.3050 0.0750 ;
        RECT 0.8850 -0.0750 1.0050 0.1800 ;
        RECT 0.5850 -0.0750 0.8850 0.0750 ;
        RECT 0.4650 -0.0750 0.5850 0.1800 ;
        RECT 0.0000 -0.0750 0.4650 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.4250 0.9750 1.4700 1.1250 ;
        RECT 1.3050 0.8175 1.4250 1.1250 ;
        RECT 1.0050 0.9750 1.3050 1.1250 ;
        RECT 0.8850 0.8625 1.0050 1.1250 ;
        RECT 0.0000 0.9750 0.8850 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.3350 0.1575 1.3950 0.2175 ;
        RECT 1.3350 0.8325 1.3950 0.8925 ;
        RECT 1.2225 0.4950 1.2825 0.5550 ;
        RECT 1.1250 0.2775 1.1850 0.3375 ;
        RECT 1.1250 0.7650 1.1850 0.8250 ;
        RECT 1.0200 0.4875 1.0800 0.5475 ;
        RECT 0.9150 0.1200 0.9750 0.1800 ;
        RECT 0.9150 0.8700 0.9750 0.9300 ;
        RECT 0.8175 0.4950 0.8775 0.5550 ;
        RECT 0.7050 0.2625 0.7650 0.3225 ;
        RECT 0.6000 0.4650 0.6600 0.5250 ;
        RECT 0.4950 0.1200 0.5550 0.1800 ;
        RECT 0.4950 0.8325 0.5550 0.8925 ;
        RECT 0.3900 0.4725 0.4500 0.5325 ;
        RECT 0.2850 0.6825 0.3450 0.7425 ;
        RECT 0.0750 0.1875 0.1350 0.2475 ;
        RECT 0.0750 0.8100 0.1350 0.8700 ;
        RECT 0.1725 0.4725 0.2325 0.5325 ;
        LAYER M1 ;
        RECT 1.0425 0.4650 1.2825 0.5850 ;
        RECT 0.9675 0.2550 1.0425 0.5850 ;
        RECT 0.7050 0.2550 0.9675 0.3375 ;
        RECT 0.8925 0.6825 0.9525 0.7875 ;
        RECT 0.8175 0.4500 0.8925 0.7875 ;
        RECT 0.7875 0.6825 0.8175 0.7875 ;
        RECT 0.6675 0.4125 0.7425 0.6000 ;
        RECT 0.3600 0.2550 0.7050 0.3300 ;
        RECT 0.5625 0.4050 0.6675 0.6000 ;
        RECT 0.2475 0.6750 0.6675 0.7500 ;
        RECT 0.1425 0.8250 0.5925 0.9000 ;
        RECT 0.3075 0.4050 0.4800 0.6000 ;
        RECT 0.2850 0.1650 0.3600 0.3300 ;
        RECT 0.0525 0.1650 0.2850 0.2700 ;
        RECT 0.0675 0.7800 0.1425 0.9000 ;
        LAYER VIA1 ;
        RECT 0.7500 0.2625 0.8250 0.3375 ;
        RECT 0.4275 0.6750 0.5025 0.7500 ;
        LAYER M2 ;
        RECT 0.5775 0.2625 0.8700 0.3375 ;
        RECT 0.5025 0.2625 0.5775 0.7500 ;
        RECT 0.3825 0.6750 0.5025 0.7500 ;
    END
END AO211_0011


MACRO AO211_0111
    CLASS CORE ;
    FOREIGN AO211_0111 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.9400 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 2.2575 0.2550 2.5725 0.7650 ;
        VIA 2.4150 0.3375 VIA12_slot ;
        VIA 2.4150 0.6825 VIA12_slot ;
        END
    END Z
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.8075 0.2625 1.9125 0.6150 ;
        RECT 1.3200 0.2625 1.8075 0.3375 ;
        RECT 1.2150 0.2625 1.3200 0.5925 ;
        VIA 1.8600 0.5325 VIA12_square ;
        VIA 1.2675 0.5175 VIA12_square ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.5450 0.4125 1.6500 0.7875 ;
        RECT 1.0500 0.7125 1.5450 0.7875 ;
        VIA 1.5975 0.5100 VIA12_square ;
        END
    END B
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.4275 0.5625 0.6675 0.6375 ;
        RECT 0.3525 0.4125 0.4275 0.6375 ;
        RECT 0.0900 0.4125 0.3525 0.4875 ;
        VIA 0.3900 0.5100 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.7875 0.2625 0.8625 0.6000 ;
        RECT 0.3525 0.2625 0.7875 0.3375 ;
        VIA 0.8250 0.5175 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 2.8875 -0.0750 2.9400 0.0750 ;
        RECT 2.7825 -0.0750 2.8875 0.3075 ;
        RECT 2.4750 -0.0750 2.7825 0.0750 ;
        RECT 2.3550 -0.0750 2.4750 0.1950 ;
        RECT 2.0475 -0.0750 2.3550 0.0750 ;
        RECT 1.9425 -0.0750 2.0475 0.2250 ;
        RECT 1.6275 -0.0750 1.9425 0.0750 ;
        RECT 1.5225 -0.0750 1.6275 0.2250 ;
        RECT 1.2150 -0.0750 1.5225 0.0750 ;
        RECT 1.0950 -0.0750 1.2150 0.2250 ;
        RECT 0.3675 -0.0750 1.0950 0.0750 ;
        RECT 0.2625 -0.0750 0.3675 0.2250 ;
        RECT 0.0000 -0.0750 0.2625 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 2.8875 0.9750 2.9400 1.1250 ;
        RECT 2.7825 0.6450 2.8875 1.1250 ;
        RECT 2.4750 0.9750 2.7825 1.1250 ;
        RECT 2.3550 0.8250 2.4750 1.1250 ;
        RECT 2.0475 0.9750 2.3550 1.1250 ;
        RECT 1.9425 0.8100 2.0475 1.1250 ;
        RECT 1.2075 0.9750 1.9425 1.1250 ;
        RECT 1.1025 0.8100 1.2075 1.1250 ;
        RECT 0.0000 0.9750 1.1025 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 2.8050 0.2175 2.8650 0.2775 ;
        RECT 2.8050 0.6675 2.8650 0.7275 ;
        RECT 2.8050 0.8325 2.8650 0.8925 ;
        RECT 2.7000 0.4800 2.7600 0.5400 ;
        RECT 2.5950 0.3075 2.6550 0.3675 ;
        RECT 2.5950 0.6525 2.6550 0.7125 ;
        RECT 2.4900 0.4800 2.5500 0.5400 ;
        RECT 2.3850 0.1275 2.4450 0.1875 ;
        RECT 2.3850 0.8325 2.4450 0.8925 ;
        RECT 2.2800 0.4800 2.3400 0.5400 ;
        RECT 2.1750 0.3075 2.2350 0.3675 ;
        RECT 2.1750 0.6525 2.2350 0.7125 ;
        RECT 2.0700 0.4800 2.1300 0.5400 ;
        RECT 1.9650 0.1425 2.0250 0.2025 ;
        RECT 1.9650 0.8325 2.0250 0.8925 ;
        RECT 1.8525 0.4950 1.9125 0.5550 ;
        RECT 1.7550 0.3075 1.8150 0.3675 ;
        RECT 1.6500 0.4800 1.7100 0.5400 ;
        RECT 1.5450 0.1425 1.6050 0.2025 ;
        RECT 1.5450 0.6600 1.6050 0.7200 ;
        RECT 1.4400 0.4800 1.5000 0.5400 ;
        RECT 1.3350 0.3075 1.3950 0.3675 ;
        RECT 1.2300 0.4800 1.2900 0.5400 ;
        RECT 1.1250 0.1575 1.1850 0.2175 ;
        RECT 1.1250 0.8325 1.1850 0.8925 ;
        RECT 0.9150 0.1725 0.9750 0.2325 ;
        RECT 0.9150 0.8175 0.9750 0.8775 ;
        RECT 0.8100 0.4950 0.8700 0.5550 ;
        RECT 0.7050 0.3000 0.7650 0.3600 ;
        RECT 0.7050 0.6750 0.7650 0.7350 ;
        RECT 0.6000 0.4875 0.6600 0.5475 ;
        RECT 0.4950 0.8325 0.5550 0.8925 ;
        RECT 0.3900 0.4800 0.4500 0.5400 ;
        RECT 0.2850 0.1425 0.3450 0.2025 ;
        RECT 0.2850 0.6600 0.3450 0.7200 ;
        RECT 0.1800 0.4800 0.2400 0.5400 ;
        RECT 0.0750 0.2925 0.1350 0.3525 ;
        RECT 0.0750 0.8175 0.1350 0.8775 ;
        LAYER M1 ;
        RECT 2.0625 0.4725 2.7900 0.5475 ;
        RECT 2.1525 0.2775 2.6850 0.3975 ;
        RECT 2.1525 0.6225 2.6850 0.7425 ;
        RECT 1.9875 0.3000 2.0625 0.5475 ;
        RECT 1.1400 0.3000 1.9875 0.3750 ;
        RECT 1.7925 0.4500 1.9125 0.7350 ;
        RECT 1.4325 0.4500 1.7175 0.5700 ;
        RECT 0.7950 0.6450 1.6500 0.7200 ;
        RECT 1.2075 0.4500 1.3575 0.5700 ;
        RECT 1.0350 0.4800 1.2075 0.5700 ;
        RECT 1.0650 0.3000 1.1400 0.4050 ;
        RECT 0.7950 0.3300 1.0650 0.4050 ;
        RECT 0.8925 0.1500 0.9975 0.2550 ;
        RECT 0.8925 0.7950 0.9975 0.9000 ;
        RECT 0.5700 0.4800 0.9300 0.5700 ;
        RECT 0.5325 0.1500 0.8925 0.2250 ;
        RECT 0.1575 0.8100 0.8925 0.9000 ;
        RECT 0.6750 0.3000 0.7950 0.4050 ;
        RECT 0.6750 0.6450 0.7950 0.7350 ;
        RECT 0.2550 0.6450 0.6750 0.7200 ;
        RECT 0.4575 0.1500 0.5325 0.3750 ;
        RECT 0.1800 0.4500 0.4650 0.5700 ;
        RECT 0.1575 0.3000 0.4575 0.3750 ;
        RECT 0.0525 0.2700 0.1575 0.3750 ;
        RECT 0.0525 0.7950 0.1575 0.9000 ;
        LAYER VIA1 ;
        RECT 2.0325 0.4725 2.1075 0.5475 ;
        RECT 0.7350 0.8100 0.8100 0.8850 ;
        LAYER M2 ;
        RECT 2.0325 0.3975 2.1075 0.9375 ;
        RECT 0.8100 0.8625 2.0325 0.9375 ;
        RECT 0.7350 0.7650 0.8100 0.9375 ;
    END
END AO211_0111


MACRO AO211_1000
    CLASS CORE ;
    FOREIGN AO211_1000 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.2600 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 1.1475 0.1500 1.2225 0.8925 ;
        RECT 1.1175 0.1500 1.1475 0.3825 ;
        RECT 1.1175 0.6675 1.1475 0.8925 ;
        END
    END Z
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.8325 0.6375 0.9075 0.9375 ;
        RECT 0.3675 0.8625 0.8325 0.9375 ;
        VIA 0.8700 0.7200 VIA12_square ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.7275 0.4125 1.1925 0.4875 ;
        RECT 0.6525 0.4125 0.7275 0.6450 ;
        VIA 0.6900 0.5175 VIA12_square ;
        END
    END B
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.4275 0.1125 0.8925 0.1875 ;
        RECT 0.3525 0.1125 0.4275 0.5250 ;
        VIA 0.3900 0.4425 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1725 0.4275 0.2325 0.5700 ;
        RECT 0.1425 0.3525 0.1725 0.5700 ;
        RECT 0.0675 0.3525 0.1425 0.6825 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.0050 -0.0750 1.2600 0.0750 ;
        RECT 0.8850 -0.0750 1.0050 0.1800 ;
        RECT 0.5850 -0.0750 0.8850 0.0750 ;
        RECT 0.4650 -0.0750 0.5850 0.1800 ;
        RECT 0.0000 -0.0750 0.4650 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.0050 0.9750 1.2600 1.1250 ;
        RECT 0.8850 0.8325 1.0050 1.1250 ;
        RECT 0.0000 0.9750 0.8850 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.1250 0.1800 1.1850 0.2400 ;
        RECT 1.1250 0.8025 1.1850 0.8625 ;
        RECT 1.0125 0.4800 1.0725 0.5400 ;
        RECT 0.9150 0.1200 0.9750 0.1800 ;
        RECT 0.9150 0.8325 0.9750 0.8925 ;
        RECT 0.8175 0.4950 0.8775 0.5550 ;
        RECT 0.7050 0.1725 0.7650 0.2325 ;
        RECT 0.6000 0.4650 0.6600 0.5250 ;
        RECT 0.4950 0.1200 0.5550 0.1800 ;
        RECT 0.4950 0.8325 0.5550 0.8925 ;
        RECT 0.3900 0.4725 0.4500 0.5325 ;
        RECT 0.1725 0.4725 0.2325 0.5325 ;
        RECT 0.0750 0.1800 0.1350 0.2400 ;
        RECT 0.0750 0.8100 0.1350 0.8700 ;
        RECT 0.2850 0.6900 0.3450 0.7500 ;
        LAYER M1 ;
        RECT 1.0425 0.4500 1.0725 0.5700 ;
        RECT 0.9675 0.2550 1.0425 0.5700 ;
        RECT 0.7875 0.2550 0.9675 0.3375 ;
        RECT 0.8925 0.6525 0.9525 0.7575 ;
        RECT 0.8175 0.4500 0.8925 0.7575 ;
        RECT 0.7875 0.6600 0.8175 0.7575 ;
        RECT 0.7050 0.1500 0.7875 0.3375 ;
        RECT 0.6675 0.4125 0.7425 0.6000 ;
        RECT 0.6825 0.1500 0.7050 0.3300 ;
        RECT 0.3600 0.2550 0.6825 0.3300 ;
        RECT 0.5625 0.4050 0.6675 0.6000 ;
        RECT 0.2475 0.6750 0.6675 0.7500 ;
        RECT 0.1425 0.8250 0.5925 0.9000 ;
        RECT 0.3075 0.4050 0.4800 0.6000 ;
        RECT 0.2850 0.1575 0.3600 0.3300 ;
        RECT 0.0525 0.1575 0.2850 0.2625 ;
        RECT 0.0675 0.7800 0.1425 0.9000 ;
        LAYER VIA1 ;
        RECT 0.7500 0.2625 0.8250 0.3375 ;
        RECT 0.4275 0.6750 0.5025 0.7500 ;
        LAYER M2 ;
        RECT 0.5775 0.2625 0.8700 0.3375 ;
        RECT 0.5025 0.2625 0.5775 0.7500 ;
        RECT 0.3825 0.6750 0.5025 0.7500 ;
    END
END AO211_1000


MACRO AO211_1010
    CLASS CORE ;
    FOREIGN AO211_1010 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.2600 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 1.1475 0.2175 1.2225 0.8325 ;
        RECT 1.1175 0.2175 1.1475 0.3825 ;
        RECT 1.1175 0.6675 1.1475 0.8325 ;
        END
    END Z
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.8325 0.6675 0.9075 0.9375 ;
        RECT 0.3675 0.8625 0.8325 0.9375 ;
        VIA 0.8700 0.7500 VIA12_square ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.7275 0.4125 1.1925 0.4875 ;
        RECT 0.6525 0.4125 0.7275 0.6450 ;
        VIA 0.6900 0.5175 VIA12_square ;
        END
    END B
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.4275 0.1125 0.8925 0.1875 ;
        RECT 0.3525 0.1125 0.4275 0.5250 ;
        VIA 0.3900 0.4425 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1725 0.4275 0.2325 0.5700 ;
        RECT 0.1425 0.3525 0.1725 0.5700 ;
        RECT 0.0675 0.3525 0.1425 0.6825 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.0050 -0.0750 1.2600 0.0750 ;
        RECT 0.8850 -0.0750 1.0050 0.1800 ;
        RECT 0.5850 -0.0750 0.8850 0.0750 ;
        RECT 0.4650 -0.0750 0.5850 0.1800 ;
        RECT 0.0000 -0.0750 0.4650 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.0050 0.9750 1.2600 1.1250 ;
        RECT 0.8850 0.8625 1.0050 1.1250 ;
        RECT 0.0000 0.9750 0.8850 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.1250 0.2700 1.1850 0.3300 ;
        RECT 1.1250 0.7200 1.1850 0.7800 ;
        RECT 1.0125 0.4800 1.0725 0.5400 ;
        RECT 0.9150 0.1200 0.9750 0.1800 ;
        RECT 0.9150 0.8700 0.9750 0.9300 ;
        RECT 0.8175 0.4950 0.8775 0.5550 ;
        RECT 0.7050 0.2625 0.7650 0.3225 ;
        RECT 0.6000 0.4650 0.6600 0.5250 ;
        RECT 0.4950 0.1200 0.5550 0.1800 ;
        RECT 0.3900 0.4725 0.4500 0.5325 ;
        RECT 0.2850 0.6825 0.3450 0.7425 ;
        RECT 0.1725 0.4725 0.2325 0.5325 ;
        RECT 0.0750 0.1875 0.1350 0.2475 ;
        RECT 0.0750 0.8100 0.1350 0.8700 ;
        RECT 0.4950 0.8325 0.5550 0.8925 ;
        LAYER M1 ;
        RECT 1.0425 0.4500 1.0725 0.5700 ;
        RECT 0.9675 0.2550 1.0425 0.5700 ;
        RECT 0.7050 0.2550 0.9675 0.3375 ;
        RECT 0.8925 0.6825 0.9525 0.7875 ;
        RECT 0.8175 0.4500 0.8925 0.7875 ;
        RECT 0.7875 0.6825 0.8175 0.7875 ;
        RECT 0.6675 0.4125 0.7425 0.6000 ;
        RECT 0.3600 0.2550 0.7050 0.3300 ;
        RECT 0.5625 0.4050 0.6675 0.6000 ;
        RECT 0.2475 0.6750 0.6675 0.7500 ;
        RECT 0.1425 0.8250 0.5925 0.9000 ;
        RECT 0.3075 0.4050 0.4800 0.6000 ;
        RECT 0.2850 0.1650 0.3600 0.3300 ;
        RECT 0.0525 0.1650 0.2850 0.2700 ;
        RECT 0.0675 0.7800 0.1425 0.9000 ;
        LAYER VIA1 ;
        RECT 0.7500 0.2625 0.8250 0.3375 ;
        RECT 0.4275 0.6750 0.5025 0.7500 ;
        LAYER M2 ;
        RECT 0.5775 0.2625 0.8700 0.3375 ;
        RECT 0.5025 0.2625 0.5775 0.7500 ;
        RECT 0.3825 0.6750 0.5025 0.7500 ;
    END
END AO211_1010


MACRO AO21_0011
    CLASS CORE ;
    FOREIGN AO21_0011 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.2600 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 1.1475 0.2925 1.2225 0.7425 ;
        RECT 0.9825 0.2925 1.1475 0.3675 ;
        RECT 0.9825 0.6675 1.1475 0.7425 ;
        RECT 0.9075 0.2175 0.9825 0.3675 ;
        RECT 0.9075 0.6675 0.9825 0.8550 ;
        END
    END Z
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.5175 0.4125 0.9825 0.4875 ;
        VIA 0.6000 0.4500 VIA12_square ;
        END
    END B
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1575 0.3675 0.2325 0.5625 ;
        RECT 0.0675 0.3675 0.1575 0.6825 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.2025 0.2625 0.6675 0.3375 ;
        VIA 0.3525 0.3000 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.2150 -0.0750 1.2600 0.0750 ;
        RECT 1.0950 -0.0750 1.2150 0.2175 ;
        RECT 0.7950 -0.0750 1.0950 0.0750 ;
        RECT 0.6750 -0.0750 0.7950 0.1800 ;
        RECT 0.1575 -0.0750 0.6750 0.0750 ;
        RECT 0.0675 -0.0750 0.1575 0.2550 ;
        RECT 0.0000 -0.0750 0.0675 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.2150 0.9750 1.2600 1.1250 ;
        RECT 1.0950 0.8175 1.2150 1.1250 ;
        RECT 0.7950 0.9750 1.0950 1.1250 ;
        RECT 0.6900 0.8250 0.7950 1.1250 ;
        RECT 0.0000 0.9750 0.6900 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.1250 0.1575 1.1850 0.2175 ;
        RECT 1.1250 0.8325 1.1850 0.8925 ;
        RECT 1.0125 0.4950 1.0725 0.5550 ;
        RECT 0.9150 0.2550 0.9750 0.3150 ;
        RECT 0.9150 0.7650 0.9750 0.8250 ;
        RECT 0.8100 0.4950 0.8700 0.5550 ;
        RECT 0.7050 0.1200 0.7650 0.1800 ;
        RECT 0.7050 0.8550 0.7650 0.9150 ;
        RECT 0.6000 0.4650 0.6600 0.5250 ;
        RECT 0.4950 0.2400 0.5550 0.3000 ;
        RECT 0.4950 0.8325 0.5550 0.8925 ;
        RECT 0.3825 0.4650 0.4425 0.5250 ;
        RECT 0.2850 0.6825 0.3450 0.7425 ;
        RECT 0.1725 0.4650 0.2325 0.5250 ;
        RECT 0.0750 0.1575 0.1350 0.2175 ;
        RECT 0.0750 0.8325 0.1350 0.8925 ;
        LAYER M1 ;
        RECT 0.8325 0.4650 1.0725 0.5850 ;
        RECT 0.7575 0.2550 0.8325 0.7500 ;
        RECT 0.5625 0.2550 0.7575 0.3300 ;
        RECT 0.3600 0.6750 0.7575 0.7500 ;
        RECT 0.5175 0.4050 0.6825 0.6000 ;
        RECT 0.1500 0.8250 0.5850 0.9000 ;
        RECT 0.4875 0.2100 0.5625 0.3300 ;
        RECT 0.3075 0.2175 0.3900 0.5700 ;
        RECT 0.2550 0.6450 0.3600 0.7500 ;
        RECT 0.0450 0.7950 0.1500 0.9000 ;
        RECT 0.3900 0.4050 0.4425 0.5700 ;
    END
END AO21_0011


MACRO AO21_0111
    CLASS CORE ;
    FOREIGN AO21_0111 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.3100 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 1.4175 0.3075 1.7325 0.7725 ;
        VIA 1.5750 0.3675 VIA12_slot ;
        VIA 1.5750 0.7125 VIA12_slot ;
        END
    END Z
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.9575 0.4125 2.2125 0.4875 ;
        RECT 1.8825 0.1125 1.9575 0.4875 ;
        RECT 1.0500 0.1125 1.8825 0.1875 ;
        RECT 0.9450 0.1125 1.0500 0.6075 ;
        VIA 2.1300 0.4500 VIA12_square ;
        VIA 0.9975 0.5250 VIA12_square ;
        END
    END B
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.5325 0.4650 0.6075 0.9375 ;
        RECT 0.0675 0.8625 0.5325 0.9375 ;
        VIA 0.5700 0.5475 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.8625 0.4500 0.8700 0.5700 ;
        RECT 0.7650 0.3450 0.8625 0.5700 ;
        RECT 0.2400 0.3450 0.7650 0.4200 ;
        RECT 0.1425 0.3450 0.2400 0.5850 ;
        RECT 0.0675 0.3450 0.1425 0.6825 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 2.0550 -0.0750 2.3100 0.0750 ;
        RECT 1.9350 -0.0750 2.0550 0.1800 ;
        RECT 1.6350 -0.0750 1.9350 0.0750 ;
        RECT 1.5150 -0.0750 1.6350 0.1875 ;
        RECT 1.2150 -0.0750 1.5150 0.0750 ;
        RECT 1.0950 -0.0750 1.2150 0.1800 ;
        RECT 0.5850 -0.0750 1.0950 0.0750 ;
        RECT 0.4650 -0.0750 0.5850 0.2700 ;
        RECT 0.0000 -0.0750 0.4650 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 2.0550 0.9750 2.3100 1.1250 ;
        RECT 1.9350 0.8700 2.0550 1.1250 ;
        RECT 1.6350 0.9750 1.9350 1.1250 ;
        RECT 1.5150 0.8550 1.6350 1.1250 ;
        RECT 1.1925 0.9750 1.5150 1.1250 ;
        RECT 1.1175 0.8400 1.1925 1.1250 ;
        RECT 0.0000 0.9750 1.1175 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 2.1750 0.2400 2.2350 0.3000 ;
        RECT 2.1750 0.7650 2.2350 0.8250 ;
        RECT 2.0700 0.4950 2.1300 0.5550 ;
        RECT 1.9650 0.1200 2.0250 0.1800 ;
        RECT 1.9650 0.8700 2.0250 0.9300 ;
        RECT 1.8600 0.4950 1.9200 0.5550 ;
        RECT 1.7550 0.2325 1.8150 0.2925 ;
        RECT 1.7550 0.7650 1.8150 0.8250 ;
        RECT 1.6500 0.4950 1.7100 0.5550 ;
        RECT 1.5450 0.1200 1.6050 0.1800 ;
        RECT 1.5450 0.8625 1.6050 0.9225 ;
        RECT 1.4400 0.4950 1.5000 0.5550 ;
        RECT 1.3350 0.2325 1.3950 0.2925 ;
        RECT 1.3350 0.7650 1.3950 0.8250 ;
        RECT 1.2300 0.4950 1.2900 0.5550 ;
        RECT 1.1250 0.1200 1.1850 0.1800 ;
        RECT 1.1250 0.8700 1.1850 0.9300 ;
        RECT 1.0200 0.4800 1.0800 0.5400 ;
        RECT 0.9150 0.1650 0.9750 0.2250 ;
        RECT 0.9150 0.8325 0.9750 0.8925 ;
        RECT 0.8100 0.4800 0.8700 0.5400 ;
        RECT 0.7050 0.6825 0.7650 0.7425 ;
        RECT 0.6000 0.4950 0.6600 0.5550 ;
        RECT 0.4950 0.1875 0.5550 0.2475 ;
        RECT 0.4950 0.8325 0.5550 0.8925 ;
        RECT 0.3900 0.4950 0.4500 0.5550 ;
        RECT 0.2850 0.6825 0.3450 0.7425 ;
        RECT 0.1800 0.4950 0.2400 0.5550 ;
        RECT 0.0750 0.1725 0.1350 0.2325 ;
        RECT 0.0750 0.8175 0.1350 0.8775 ;
        LAYER M1 ;
        RECT 2.1675 0.2100 2.2425 0.3300 ;
        RECT 2.0475 0.4050 2.2425 0.6150 ;
        RECT 2.1675 0.6900 2.2425 0.8625 ;
        RECT 1.9725 0.2550 2.1675 0.3300 ;
        RECT 1.8975 0.6900 2.1675 0.7950 ;
        RECT 1.8975 0.2550 1.9725 0.5700 ;
        RECT 1.2300 0.4950 1.8975 0.5700 ;
        RECT 1.7475 0.1800 1.8225 0.4200 ;
        RECT 1.7475 0.6675 1.8225 0.8550 ;
        RECT 1.4025 0.3075 1.7475 0.4200 ;
        RECT 1.4175 0.6675 1.7475 0.7575 ;
        RECT 1.3125 0.6675 1.4175 0.8550 ;
        RECT 1.3275 0.1800 1.4025 0.4200 ;
        RECT 1.1550 0.2550 1.2300 0.5700 ;
        RECT 1.0200 0.2550 1.1550 0.3300 ;
        RECT 0.9450 0.4050 1.0800 0.6600 ;
        RECT 0.9300 0.7350 1.0425 0.9000 ;
        RECT 0.9450 0.1500 1.0200 0.3300 ;
        RECT 0.6825 0.1500 0.9450 0.2550 ;
        RECT 0.1575 0.8250 0.9300 0.9000 ;
        RECT 0.2475 0.6750 0.8175 0.7500 ;
        RECT 0.3600 0.4950 0.6900 0.6000 ;
        RECT 0.0525 0.1500 0.3675 0.2550 ;
        RECT 0.0525 0.7950 0.1575 0.9000 ;
        LAYER VIA1 ;
        RECT 1.9425 0.7125 2.0175 0.7875 ;
        RECT 0.9375 0.7800 1.0125 0.8550 ;
        RECT 0.7275 0.1800 0.8025 0.2550 ;
        RECT 0.6975 0.6750 0.7725 0.7500 ;
        RECT 0.2475 0.1800 0.3225 0.2550 ;
        LAYER M2 ;
        RECT 1.9425 0.7125 2.0625 0.7875 ;
        RECT 1.8600 0.7125 1.9425 0.9375 ;
        RECT 1.0275 0.8625 1.8600 0.9375 ;
        RECT 0.9225 0.7350 1.0275 0.9375 ;
        RECT 0.7875 0.1650 0.8475 0.2700 ;
        RECT 0.6825 0.1650 0.7875 0.7875 ;
        RECT 0.1800 0.1650 0.6825 0.2550 ;
    END
END AO21_0111


MACRO AO21_1000
    CLASS CORE ;
    FOREIGN AO21_1000 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.0500 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.9375 0.1500 1.0125 0.9000 ;
        RECT 0.9075 0.1500 0.9375 0.3825 ;
        RECT 0.9075 0.6675 0.9375 0.9000 ;
        END
    END Z
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.5175 0.4125 0.9825 0.4875 ;
        VIA 0.6000 0.4500 VIA12_square ;
        END
    END B
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1575 0.3675 0.2325 0.5625 ;
        RECT 0.0675 0.3675 0.1575 0.6825 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.2025 0.2625 0.6675 0.3375 ;
        VIA 0.3525 0.3000 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.7950 -0.0750 1.0500 0.0750 ;
        RECT 0.6750 -0.0750 0.7950 0.1800 ;
        RECT 0.1575 -0.0750 0.6750 0.0750 ;
        RECT 0.0675 -0.0750 0.1575 0.2550 ;
        RECT 0.0000 -0.0750 0.0675 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.7950 0.9750 1.0500 1.1250 ;
        RECT 0.6900 0.8250 0.7950 1.1250 ;
        RECT 0.0000 0.9750 0.6900 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 0.9150 0.1800 0.9750 0.2400 ;
        RECT 0.9150 0.8025 0.9750 0.8625 ;
        RECT 0.8025 0.4875 0.8625 0.5475 ;
        RECT 0.7050 0.1200 0.7650 0.1800 ;
        RECT 0.7050 0.8550 0.7650 0.9150 ;
        RECT 0.6000 0.4650 0.6600 0.5250 ;
        RECT 0.4950 0.1800 0.5550 0.2400 ;
        RECT 0.4950 0.8250 0.5550 0.8850 ;
        RECT 0.3825 0.4650 0.4425 0.5250 ;
        RECT 0.2850 0.6900 0.3450 0.7500 ;
        RECT 0.1725 0.4650 0.2325 0.5250 ;
        RECT 0.0750 0.1575 0.1350 0.2175 ;
        RECT 0.0750 0.8175 0.1350 0.8775 ;
        LAYER M1 ;
        RECT 0.8325 0.4575 0.8625 0.5775 ;
        RECT 0.5775 0.2550 0.7575 0.3300 ;
        RECT 0.3600 0.6750 0.7575 0.7500 ;
        RECT 0.5175 0.4050 0.6825 0.6000 ;
        RECT 0.1575 0.8250 0.5850 0.9000 ;
        RECT 0.4725 0.1500 0.5775 0.3300 ;
        RECT 0.3900 0.4050 0.4425 0.5700 ;
        RECT 0.3075 0.2175 0.3900 0.5700 ;
        RECT 0.2550 0.6450 0.3600 0.7500 ;
        RECT 0.0525 0.7950 0.1575 0.9000 ;
        RECT 0.7575 0.2550 0.8325 0.7500 ;
    END
END AO21_1000


MACRO AO21_1010
    CLASS CORE ;
    FOREIGN AO21_1010 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.0500 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.9375 0.2175 1.0125 0.8325 ;
        RECT 0.9075 0.2175 0.9375 0.3825 ;
        RECT 0.9075 0.6675 0.9375 0.8325 ;
        END
    END Z
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.5175 0.4125 0.9825 0.4875 ;
        VIA 0.6000 0.4500 VIA12_square ;
        END
    END B
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1575 0.3675 0.2325 0.5625 ;
        RECT 0.0675 0.3675 0.1575 0.6825 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.2025 0.2625 0.6675 0.3375 ;
        VIA 0.3525 0.3000 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.7950 -0.0750 1.0500 0.0750 ;
        RECT 0.6750 -0.0750 0.7950 0.1800 ;
        RECT 0.1575 -0.0750 0.6750 0.0750 ;
        RECT 0.0675 -0.0750 0.1575 0.2550 ;
        RECT 0.0000 -0.0750 0.0675 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.7950 0.9750 1.0500 1.1250 ;
        RECT 0.6900 0.8250 0.7950 1.1250 ;
        RECT 0.0000 0.9750 0.6900 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 0.9150 0.2700 0.9750 0.3300 ;
        RECT 0.9150 0.7200 0.9750 0.7800 ;
        RECT 0.8025 0.4875 0.8625 0.5475 ;
        RECT 0.7050 0.1200 0.7650 0.1800 ;
        RECT 0.7050 0.8550 0.7650 0.9150 ;
        RECT 0.6000 0.4650 0.6600 0.5250 ;
        RECT 0.4950 0.2400 0.5550 0.3000 ;
        RECT 0.4950 0.8325 0.5550 0.8925 ;
        RECT 0.3825 0.4650 0.4425 0.5250 ;
        RECT 0.2850 0.6825 0.3450 0.7425 ;
        RECT 0.1725 0.4650 0.2325 0.5250 ;
        RECT 0.0750 0.1575 0.1350 0.2175 ;
        RECT 0.0750 0.8325 0.1350 0.8925 ;
        LAYER M1 ;
        RECT 0.8325 0.4575 0.8625 0.5775 ;
        RECT 0.5625 0.2550 0.7575 0.3300 ;
        RECT 0.3600 0.6750 0.7575 0.7500 ;
        RECT 0.5175 0.4050 0.6825 0.6000 ;
        RECT 0.1500 0.8250 0.5850 0.9000 ;
        RECT 0.4875 0.2100 0.5625 0.3300 ;
        RECT 0.3900 0.4050 0.4425 0.5700 ;
        RECT 0.3075 0.2175 0.3900 0.5700 ;
        RECT 0.2550 0.6450 0.3600 0.7500 ;
        RECT 0.0450 0.7950 0.1500 0.9000 ;
        RECT 0.7575 0.2550 0.8325 0.7500 ;
    END
END AO21_1010


MACRO AO221_0011
    CLASS CORE ;
    FOREIGN AO221_0011 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.8900 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 1.7775 0.3075 1.8525 0.7425 ;
        RECT 1.6125 0.3075 1.7775 0.3825 ;
        RECT 1.6125 0.6675 1.7775 0.7425 ;
        RECT 1.5375 0.2175 1.6125 0.3825 ;
        RECT 1.5375 0.6675 1.6125 0.8325 ;
        END
    END Z
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.1475 0.1125 1.6125 0.1875 ;
        RECT 1.0725 0.1125 1.1475 0.4500 ;
        RECT 0.7275 0.3750 1.0725 0.4500 ;
        RECT 0.6525 0.3750 0.7275 0.5625 ;
        VIA 0.6900 0.4800 VIA12_square ;
        END
    END C
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.8775 0.8625 1.4175 0.9375 ;
        RECT 0.8775 0.5250 0.9675 0.6300 ;
        RECT 0.8025 0.5250 0.8775 0.9375 ;
        VIA 0.8850 0.5775 VIA12_square ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.1475 0.7125 1.6125 0.7875 ;
        RECT 1.1475 0.5625 1.2825 0.6375 ;
        RECT 1.0725 0.5625 1.1475 0.7875 ;
        VIA 1.1850 0.6000 VIA12_square ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1425 0.4425 0.2475 0.5625 ;
        RECT 0.0675 0.3675 0.1425 0.6825 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.4275 0.8625 0.6075 0.9375 ;
        RECT 0.3525 0.3900 0.4275 0.9375 ;
        RECT 0.0675 0.8625 0.3525 0.9375 ;
        VIA 0.3900 0.4725 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.8450 -0.0750 1.8900 0.0750 ;
        RECT 1.7250 -0.0750 1.8450 0.2175 ;
        RECT 1.4250 -0.0750 1.7250 0.0750 ;
        RECT 1.3050 -0.0750 1.4250 0.2175 ;
        RECT 0.7650 -0.0750 1.3050 0.0750 ;
        RECT 0.6600 -0.0750 0.7650 0.2400 ;
        RECT 0.1650 -0.0750 0.6600 0.0750 ;
        RECT 0.0450 -0.0750 0.1650 0.2325 ;
        RECT 0.0000 -0.0750 0.0450 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.8450 0.9750 1.8900 1.1250 ;
        RECT 1.7250 0.8325 1.8450 1.1250 ;
        RECT 1.4250 0.9750 1.7250 1.1250 ;
        RECT 1.3050 0.7275 1.4250 1.1250 ;
        RECT 1.0050 0.9750 1.3050 1.1250 ;
        RECT 0.8850 0.8700 1.0050 1.1250 ;
        RECT 0.0000 0.9750 0.8850 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.7550 0.1575 1.8150 0.2175 ;
        RECT 1.7550 0.8325 1.8150 0.8925 ;
        RECT 1.6425 0.4875 1.7025 0.5475 ;
        RECT 1.5450 0.2700 1.6050 0.3300 ;
        RECT 1.5450 0.7200 1.6050 0.7800 ;
        RECT 1.4400 0.4875 1.5000 0.5475 ;
        RECT 1.3350 0.1575 1.3950 0.2175 ;
        RECT 1.3350 0.7575 1.3950 0.8175 ;
        RECT 1.1250 0.2175 1.1850 0.2775 ;
        RECT 1.1250 0.7575 1.1850 0.8175 ;
        RECT 1.0275 0.4950 1.0875 0.5550 ;
        RECT 0.9150 0.8700 0.9750 0.9300 ;
        RECT 0.8100 0.4875 0.8700 0.5475 ;
        RECT 0.7050 0.1500 0.7650 0.2100 ;
        RECT 0.7050 0.7575 0.7650 0.8175 ;
        RECT 0.6000 0.4650 0.6600 0.5250 ;
        RECT 0.4950 0.1800 0.5550 0.2400 ;
        RECT 0.4950 0.8325 0.5550 0.8925 ;
        RECT 0.3900 0.4650 0.4500 0.5250 ;
        RECT 0.2850 0.6525 0.3450 0.7125 ;
        RECT 0.1800 0.4725 0.2400 0.5325 ;
        RECT 0.0750 0.1575 0.1350 0.2175 ;
        RECT 0.0750 0.8250 0.1350 0.8850 ;
        LAYER M1 ;
        RECT 1.4625 0.4575 1.7025 0.5775 ;
        RECT 1.3875 0.2925 1.4625 0.5775 ;
        RECT 1.1925 0.2925 1.3875 0.3675 ;
        RECT 1.1325 0.5325 1.2825 0.6375 ;
        RECT 1.1175 0.1575 1.1925 0.3675 ;
        RECT 1.0950 0.7200 1.1850 0.8550 ;
        RECT 1.0275 0.4500 1.1325 0.6375 ;
        RECT 0.8400 0.1575 1.1175 0.2625 ;
        RECT 0.7950 0.7200 1.0950 0.7950 ;
        RECT 0.8100 0.3525 0.9525 0.6450 ;
        RECT 0.6975 0.7200 0.7950 0.8475 ;
        RECT 0.5775 0.3450 0.7350 0.5625 ;
        RECT 0.3825 0.6375 0.6225 0.7500 ;
        RECT 0.2775 0.1575 0.5850 0.2700 ;
        RECT 0.1500 0.8250 0.5850 0.9000 ;
        RECT 0.3375 0.3450 0.5025 0.5550 ;
        RECT 0.2400 0.6450 0.3825 0.7500 ;
        RECT 0.0450 0.7950 0.1500 0.9000 ;
        LAYER VIA1 ;
        RECT 0.8850 0.1875 0.9600 0.2625 ;
        RECT 0.5025 0.6375 0.5775 0.7125 ;
        RECT 0.4275 0.1575 0.5025 0.2325 ;
        LAYER M2 ;
        RECT 0.8400 0.1575 0.9900 0.3000 ;
        RECT 0.5775 0.2250 0.8400 0.3000 ;
        RECT 0.5775 0.7125 0.6075 0.7875 ;
        RECT 0.5025 0.1575 0.5775 0.7875 ;
        RECT 0.3825 0.1575 0.5025 0.2325 ;
    END
END AO221_0011


MACRO AO221_0111
    CLASS CORE ;
    FOREIGN AO221_0111 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.3600 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 2.6775 0.2400 2.9925 0.7500 ;
        VIA 2.8350 0.3225 VIA12_slot ;
        VIA 2.8350 0.6675 VIA12_slot ;
        END
    END Z
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.1025 0.4275 1.2075 0.9375 ;
        RECT 0.6375 0.8625 1.1025 0.9375 ;
        VIA 1.1550 0.5250 VIA12_square ;
        END
    END C
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.6275 0.8625 2.0925 0.9375 ;
        RECT 1.5225 0.3600 1.6275 0.9375 ;
        VIA 1.5750 0.4725 VIA12_square ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 2.0475 0.7125 2.5125 0.7875 ;
        RECT 1.9425 0.4200 2.0475 0.7875 ;
        VIA 1.9950 0.5250 VIA12_square ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.8025 0.3450 0.8775 0.5700 ;
        RECT 0.2400 0.3450 0.8025 0.4200 ;
        RECT 0.1425 0.3450 0.2400 0.5550 ;
        RECT 0.0675 0.3450 0.1425 0.6825 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.4875 0.4650 0.5625 0.7875 ;
        RECT 0.0975 0.7125 0.4875 0.7875 ;
        VIA 0.5250 0.5475 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 3.2925 -0.0750 3.3600 0.0750 ;
        RECT 3.2175 -0.0750 3.2925 0.3150 ;
        RECT 2.8950 -0.0750 3.2175 0.0750 ;
        RECT 2.7750 -0.0750 2.8950 0.1950 ;
        RECT 2.4750 -0.0750 2.7750 0.0750 ;
        RECT 2.3550 -0.0750 2.4750 0.2475 ;
        RECT 1.6350 -0.0750 2.3550 0.0750 ;
        RECT 1.5150 -0.0750 1.6350 0.2475 ;
        RECT 1.4100 -0.0750 1.5150 0.0750 ;
        RECT 1.3200 -0.0750 1.4100 0.3075 ;
        RECT 1.0200 -0.0750 1.3200 0.0750 ;
        RECT 0.9150 -0.0750 1.0200 0.2550 ;
        RECT 0.1575 -0.0750 0.9150 0.0750 ;
        RECT 0.0525 -0.0750 0.1575 0.2475 ;
        RECT 0.0000 -0.0750 0.0525 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 3.2925 0.9750 3.3600 1.1250 ;
        RECT 3.2175 0.6375 3.2925 1.1250 ;
        RECT 2.8725 0.9750 3.2175 1.1250 ;
        RECT 2.7975 0.8175 2.8725 1.1250 ;
        RECT 2.4525 0.9750 2.7975 1.1250 ;
        RECT 2.3775 0.6375 2.4525 1.1250 ;
        RECT 2.0550 0.9750 2.3775 1.1250 ;
        RECT 1.9350 0.8025 2.0550 1.1250 ;
        RECT 1.6350 0.9750 1.9350 1.1250 ;
        RECT 1.5300 0.8025 1.6350 1.1250 ;
        RECT 0.0000 0.9750 1.5300 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 3.2250 0.2250 3.2850 0.2850 ;
        RECT 3.2250 0.6675 3.2850 0.7275 ;
        RECT 3.2250 0.8325 3.2850 0.8925 ;
        RECT 3.1200 0.4650 3.1800 0.5250 ;
        RECT 3.0150 0.2250 3.0750 0.2850 ;
        RECT 3.0150 0.7575 3.0750 0.8175 ;
        RECT 2.9100 0.4650 2.9700 0.5250 ;
        RECT 2.8050 0.1275 2.8650 0.1875 ;
        RECT 2.8050 0.8475 2.8650 0.9075 ;
        RECT 2.7000 0.4650 2.7600 0.5250 ;
        RECT 2.5950 0.2250 2.6550 0.2850 ;
        RECT 2.5950 0.7575 2.6550 0.8175 ;
        RECT 2.4900 0.4650 2.5500 0.5250 ;
        RECT 2.3850 0.1650 2.4450 0.2250 ;
        RECT 2.3850 0.6675 2.4450 0.7275 ;
        RECT 2.3850 0.8325 2.4450 0.8925 ;
        RECT 2.2800 0.4650 2.3400 0.5250 ;
        RECT 2.1750 0.6675 2.2350 0.7275 ;
        RECT 2.0700 0.4950 2.1300 0.5550 ;
        RECT 1.9650 0.1725 2.0250 0.2325 ;
        RECT 1.9650 0.8325 2.0250 0.8925 ;
        RECT 1.8600 0.4875 1.9200 0.5475 ;
        RECT 1.7550 0.6600 1.8150 0.7200 ;
        RECT 1.6500 0.4650 1.7100 0.5250 ;
        RECT 1.5450 0.1725 1.6050 0.2325 ;
        RECT 1.5450 0.8325 1.6050 0.8925 ;
        RECT 1.3350 0.2025 1.3950 0.2625 ;
        RECT 1.3350 0.8325 1.3950 0.8925 ;
        RECT 1.2300 0.4875 1.2900 0.5475 ;
        RECT 1.1250 0.1800 1.1850 0.2400 ;
        RECT 1.1250 0.6600 1.1850 0.7200 ;
        RECT 1.0200 0.4875 1.0800 0.5475 ;
        RECT 0.9150 0.1650 0.9750 0.2250 ;
        RECT 0.9150 0.8325 0.9750 0.8925 ;
        RECT 0.8100 0.4800 0.8700 0.5400 ;
        RECT 0.7050 0.6825 0.7650 0.7425 ;
        RECT 0.6000 0.4950 0.6600 0.5550 ;
        RECT 0.4950 0.1875 0.5550 0.2475 ;
        RECT 0.4950 0.8325 0.5550 0.8925 ;
        RECT 0.3900 0.4950 0.4500 0.5550 ;
        RECT 0.2850 0.6825 0.3450 0.7425 ;
        RECT 0.1800 0.4650 0.2400 0.5250 ;
        RECT 0.0750 0.1575 0.1350 0.2175 ;
        RECT 0.0750 0.8175 0.1350 0.8775 ;
        LAYER M1 ;
        RECT 2.4900 0.4425 3.2100 0.5475 ;
        RECT 2.9925 0.1950 3.0975 0.3675 ;
        RECT 3.0075 0.6225 3.0825 0.8700 ;
        RECT 2.6625 0.6225 3.0075 0.7125 ;
        RECT 2.6775 0.2775 2.9925 0.3675 ;
        RECT 2.5725 0.1950 2.6775 0.3675 ;
        RECT 2.5875 0.6225 2.6625 0.8700 ;
        RECT 2.4150 0.3750 2.4900 0.5475 ;
        RECT 2.2350 0.3225 2.3400 0.5550 ;
        RECT 1.0950 0.6525 2.2650 0.7275 ;
        RECT 1.7100 0.3225 2.2350 0.3975 ;
        RECT 1.8225 0.1500 2.1675 0.2475 ;
        RECT 1.8300 0.4725 2.1525 0.5775 ;
        RECT 1.6350 0.3225 1.7100 0.5550 ;
        RECT 1.5375 0.3900 1.6350 0.5550 ;
        RECT 0.1575 0.8250 1.4250 0.9000 ;
        RECT 0.9900 0.4800 1.3200 0.5775 ;
        RECT 1.0950 0.1650 1.2450 0.3975 ;
        RECT 0.2475 0.6750 0.8550 0.7500 ;
        RECT 0.4650 0.1650 0.8400 0.2700 ;
        RECT 0.3600 0.4950 0.6900 0.6000 ;
        RECT 0.0525 0.7950 0.1575 0.9000 ;
        LAYER VIA1 ;
        RECT 2.4150 0.4275 2.4900 0.5025 ;
        RECT 1.9575 0.1650 2.0325 0.2400 ;
        RECT 1.1325 0.1800 1.2075 0.2550 ;
        RECT 0.7350 0.6750 0.8100 0.7500 ;
        RECT 0.7275 0.1800 0.8025 0.2550 ;
        LAYER M2 ;
        RECT 2.3775 0.1650 2.5050 0.5400 ;
        RECT 0.7800 0.1650 2.3775 0.2700 ;
        RECT 0.7800 0.6750 0.8550 0.7500 ;
        RECT 0.6900 0.1650 0.7800 0.7500 ;
    END
END AO221_0111


MACRO AO221_1000
    CLASS CORE ;
    FOREIGN AO221_1000 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.6800 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 1.5675 0.1500 1.6425 0.9000 ;
        RECT 1.5375 0.1500 1.5675 0.3825 ;
        RECT 1.5375 0.6675 1.5675 0.9000 ;
        END
    END Z
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.1475 0.1125 1.6125 0.1875 ;
        RECT 1.0725 0.1125 1.1475 0.4500 ;
        RECT 0.7275 0.3750 1.0725 0.4500 ;
        RECT 0.6525 0.3750 0.7275 0.5625 ;
        VIA 0.6900 0.4800 VIA12_square ;
        END
    END C
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.8775 0.8625 1.4175 0.9375 ;
        RECT 0.8775 0.5250 0.9675 0.6300 ;
        RECT 0.8025 0.5250 0.8775 0.9375 ;
        VIA 0.8850 0.5775 VIA12_square ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.1475 0.7125 1.6125 0.7875 ;
        RECT 1.1475 0.5625 1.2825 0.6375 ;
        RECT 1.0725 0.5625 1.1475 0.7875 ;
        VIA 1.1850 0.6000 VIA12_square ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1425 0.4425 0.2475 0.5625 ;
        RECT 0.0675 0.3675 0.1425 0.6825 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.4275 0.8625 0.6075 0.9375 ;
        RECT 0.3525 0.3900 0.4275 0.9375 ;
        RECT 0.0675 0.8625 0.3525 0.9375 ;
        VIA 0.3900 0.4725 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.4250 -0.0750 1.6800 0.0750 ;
        RECT 1.3050 -0.0750 1.4250 0.2175 ;
        RECT 0.7650 -0.0750 1.3050 0.0750 ;
        RECT 0.6600 -0.0750 0.7650 0.2400 ;
        RECT 0.1650 -0.0750 0.6600 0.0750 ;
        RECT 0.0450 -0.0750 0.1650 0.2325 ;
        RECT 0.0000 -0.0750 0.0450 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.4250 0.9750 1.6800 1.1250 ;
        RECT 1.3050 0.7275 1.4250 1.1250 ;
        RECT 1.0050 0.9750 1.3050 1.1250 ;
        RECT 0.8850 0.8700 1.0050 1.1250 ;
        RECT 0.0000 0.9750 0.8850 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.5450 0.1800 1.6050 0.2400 ;
        RECT 1.5450 0.8100 1.6050 0.8700 ;
        RECT 1.4325 0.4725 1.4925 0.5325 ;
        RECT 1.3350 0.1575 1.3950 0.2175 ;
        RECT 1.3350 0.8100 1.3950 0.8700 ;
        RECT 1.1250 0.1800 1.1850 0.2400 ;
        RECT 1.1250 0.8100 1.1850 0.8700 ;
        RECT 1.0275 0.4950 1.0875 0.5550 ;
        RECT 0.9150 0.8700 0.9750 0.9300 ;
        RECT 0.8100 0.4875 0.8700 0.5475 ;
        RECT 0.7050 0.1500 0.7650 0.2100 ;
        RECT 0.7050 0.8025 0.7650 0.8625 ;
        RECT 0.6000 0.4650 0.6600 0.5250 ;
        RECT 0.4950 0.1800 0.5550 0.2400 ;
        RECT 0.4950 0.8325 0.5550 0.8925 ;
        RECT 0.3900 0.4650 0.4500 0.5250 ;
        RECT 0.2850 0.6825 0.3450 0.7425 ;
        RECT 0.1800 0.4725 0.2400 0.5325 ;
        RECT 0.0750 0.1575 0.1350 0.2175 ;
        RECT 0.0750 0.8250 0.1350 0.8850 ;
        LAYER M1 ;
        RECT 1.4625 0.4425 1.4925 0.5625 ;
        RECT 1.3875 0.2925 1.4625 0.5625 ;
        RECT 1.1925 0.2925 1.3875 0.3675 ;
        RECT 1.1325 0.5325 1.2825 0.6375 ;
        RECT 1.1175 0.1500 1.1925 0.3675 ;
        RECT 1.0800 0.7200 1.1850 0.9000 ;
        RECT 1.0275 0.4500 1.1325 0.6375 ;
        RECT 0.8400 0.1500 1.1175 0.2625 ;
        RECT 0.8025 0.7200 1.0800 0.7950 ;
        RECT 0.8100 0.3525 0.9525 0.6450 ;
        RECT 0.6975 0.7200 0.8025 0.8925 ;
        RECT 0.5775 0.3450 0.7350 0.5625 ;
        RECT 0.3825 0.6375 0.6225 0.7500 ;
        RECT 0.2775 0.1575 0.5850 0.2700 ;
        RECT 0.1500 0.8250 0.5850 0.9000 ;
        RECT 0.3375 0.3450 0.5025 0.5550 ;
        RECT 0.2400 0.6450 0.3825 0.7500 ;
        RECT 0.0450 0.7950 0.1500 0.9000 ;
        LAYER VIA1 ;
        RECT 0.8850 0.1875 0.9600 0.2625 ;
        RECT 0.5025 0.6375 0.5775 0.7125 ;
        RECT 0.4275 0.1575 0.5025 0.2325 ;
        LAYER M2 ;
        RECT 0.8400 0.1575 0.9900 0.3000 ;
        RECT 0.5775 0.2250 0.8400 0.3000 ;
        RECT 0.5775 0.7125 0.6075 0.7875 ;
        RECT 0.5025 0.1575 0.5775 0.7875 ;
        RECT 0.3825 0.1575 0.5025 0.2325 ;
    END
END AO221_1000


MACRO AO221_1010
    CLASS CORE ;
    FOREIGN AO221_1010 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.6800 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 1.5675 0.2175 1.6425 0.8325 ;
        RECT 1.5375 0.2175 1.5675 0.3825 ;
        RECT 1.5375 0.6675 1.5675 0.8325 ;
        END
    END Z
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.1475 0.1125 1.6125 0.1875 ;
        RECT 1.0725 0.1125 1.1475 0.4500 ;
        RECT 0.7275 0.3750 1.0725 0.4500 ;
        RECT 0.6525 0.3750 0.7275 0.5625 ;
        VIA 0.6900 0.4800 VIA12_square ;
        END
    END C
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.8775 0.8625 1.4175 0.9375 ;
        RECT 0.8775 0.5250 0.9675 0.6300 ;
        RECT 0.8025 0.5250 0.8775 0.9375 ;
        VIA 0.8850 0.5775 VIA12_square ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.1475 0.7125 1.6125 0.7875 ;
        RECT 1.1475 0.5625 1.2825 0.6375 ;
        RECT 1.0725 0.5625 1.1475 0.7875 ;
        VIA 1.1850 0.6000 VIA12_square ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1425 0.4425 0.2475 0.5625 ;
        RECT 0.0675 0.3675 0.1425 0.6825 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.4275 0.8625 0.6075 0.9375 ;
        RECT 0.3525 0.3900 0.4275 0.9375 ;
        RECT 0.0675 0.8625 0.3525 0.9375 ;
        VIA 0.3900 0.4725 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.4250 -0.0750 1.6800 0.0750 ;
        RECT 1.3050 -0.0750 1.4250 0.2175 ;
        RECT 0.7650 -0.0750 1.3050 0.0750 ;
        RECT 0.6600 -0.0750 0.7650 0.2400 ;
        RECT 0.1650 -0.0750 0.6600 0.0750 ;
        RECT 0.0450 -0.0750 0.1650 0.2325 ;
        RECT 0.0000 -0.0750 0.0450 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.4250 0.9750 1.6800 1.1250 ;
        RECT 1.3050 0.7275 1.4250 1.1250 ;
        RECT 1.0050 0.9750 1.3050 1.1250 ;
        RECT 0.8850 0.8700 1.0050 1.1250 ;
        RECT 0.0000 0.9750 0.8850 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.5450 0.2700 1.6050 0.3300 ;
        RECT 1.5450 0.7200 1.6050 0.7800 ;
        RECT 1.4325 0.4725 1.4925 0.5325 ;
        RECT 1.3350 0.1575 1.3950 0.2175 ;
        RECT 1.3350 0.7575 1.3950 0.8175 ;
        RECT 1.1250 0.2175 1.1850 0.2775 ;
        RECT 1.1250 0.7575 1.1850 0.8175 ;
        RECT 1.0275 0.4950 1.0875 0.5550 ;
        RECT 0.9150 0.8700 0.9750 0.9300 ;
        RECT 0.8100 0.4875 0.8700 0.5475 ;
        RECT 0.7050 0.1500 0.7650 0.2100 ;
        RECT 0.7050 0.7575 0.7650 0.8175 ;
        RECT 0.6000 0.4650 0.6600 0.5250 ;
        RECT 0.4950 0.1800 0.5550 0.2400 ;
        RECT 0.4950 0.8325 0.5550 0.8925 ;
        RECT 0.3900 0.4650 0.4500 0.5250 ;
        RECT 0.2850 0.6525 0.3450 0.7125 ;
        RECT 0.1800 0.4725 0.2400 0.5325 ;
        RECT 0.0750 0.1575 0.1350 0.2175 ;
        RECT 0.0750 0.8250 0.1350 0.8850 ;
        LAYER M1 ;
        RECT 1.4625 0.4425 1.4925 0.5625 ;
        RECT 1.3875 0.2925 1.4625 0.5625 ;
        RECT 1.1925 0.2925 1.3875 0.3675 ;
        RECT 1.1325 0.5325 1.2825 0.6375 ;
        RECT 1.1175 0.1575 1.1925 0.3675 ;
        RECT 1.0950 0.7200 1.1850 0.8550 ;
        RECT 1.0275 0.4500 1.1325 0.6375 ;
        RECT 0.8400 0.1575 1.1175 0.2625 ;
        RECT 0.7950 0.7200 1.0950 0.7950 ;
        RECT 0.8100 0.3525 0.9525 0.6450 ;
        RECT 0.6975 0.7200 0.7950 0.8475 ;
        RECT 0.5775 0.3450 0.7350 0.5625 ;
        RECT 0.3825 0.6375 0.6225 0.7500 ;
        RECT 0.2775 0.1575 0.5850 0.2700 ;
        RECT 0.1500 0.8250 0.5850 0.9000 ;
        RECT 0.3375 0.3450 0.5025 0.5550 ;
        RECT 0.2400 0.6450 0.3825 0.7500 ;
        RECT 0.0450 0.7950 0.1500 0.9000 ;
        LAYER VIA1 ;
        RECT 0.8850 0.1875 0.9600 0.2625 ;
        RECT 0.5025 0.6375 0.5775 0.7125 ;
        RECT 0.4275 0.1575 0.5025 0.2325 ;
        LAYER M2 ;
        RECT 0.8400 0.1575 0.9900 0.3000 ;
        RECT 0.5775 0.2250 0.8400 0.3000 ;
        RECT 0.5775 0.7125 0.6075 0.7875 ;
        RECT 0.5025 0.1575 0.5775 0.7875 ;
        RECT 0.3825 0.1575 0.5025 0.2325 ;
    END
END AO221_1010


MACRO AO222_0011
    CLASS CORE ;
    FOREIGN AO222_0011 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.1000 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 1.9875 0.3075 2.0625 0.7425 ;
        RECT 1.8225 0.3075 1.9875 0.3825 ;
        RECT 1.8225 0.6675 1.9875 0.7425 ;
        RECT 1.7475 0.2175 1.8225 0.3825 ;
        RECT 1.7475 0.6675 1.8225 0.8550 ;
        END
    END Z
    PIN C2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.2000 0.5625 1.6650 0.6375 ;
        VIA 1.4625 0.6000 VIA12_square ;
        END
    END C2
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.0575 0.4125 1.5225 0.4875 ;
        VIA 1.1700 0.4500 VIA12_square ;
        END
    END C1
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.9375 0.7125 1.4025 0.7875 ;
        RECT 0.8625 0.4050 0.9375 0.7875 ;
        VIA 0.9000 0.4875 VIA12_square ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.6150 0.3600 0.6375 0.5100 ;
        RECT 0.5325 0.1125 0.6150 0.5100 ;
        RECT 0.0675 0.1125 0.5325 0.1875 ;
        VIA 0.5850 0.4350 VIA12_square ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1425 0.4350 0.2325 0.5550 ;
        RECT 0.0675 0.3675 0.1425 0.6825 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.4275 0.8625 0.8925 0.9375 ;
        RECT 0.3525 0.4050 0.4275 0.9375 ;
        VIA 0.3900 0.4875 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 2.0550 -0.0750 2.1000 0.0750 ;
        RECT 1.9350 -0.0750 2.0550 0.2175 ;
        RECT 1.6350 -0.0750 1.9350 0.0750 ;
        RECT 1.5150 -0.0750 1.6350 0.1800 ;
        RECT 0.9975 -0.0750 1.5150 0.0750 ;
        RECT 0.8925 -0.0750 0.9975 0.2400 ;
        RECT 0.1425 -0.0750 0.8925 0.0750 ;
        RECT 0.0675 -0.0750 0.1425 0.2625 ;
        RECT 0.0000 -0.0750 0.0675 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 2.0550 0.9750 2.1000 1.1250 ;
        RECT 1.9350 0.8175 2.0550 1.1250 ;
        RECT 1.6350 0.9750 1.9350 1.1250 ;
        RECT 1.5150 0.8250 1.6350 1.1250 ;
        RECT 1.1850 0.9750 1.5150 1.1250 ;
        RECT 1.0800 0.8025 1.1850 1.1250 ;
        RECT 0.0000 0.9750 1.0800 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.9650 0.1575 2.0250 0.2175 ;
        RECT 1.9650 0.8325 2.0250 0.8925 ;
        RECT 1.8525 0.4950 1.9125 0.5550 ;
        RECT 1.7550 0.2550 1.8150 0.3150 ;
        RECT 1.7550 0.7650 1.8150 0.8250 ;
        RECT 1.6500 0.4950 1.7100 0.5550 ;
        RECT 1.5450 0.1200 1.6050 0.1800 ;
        RECT 1.5450 0.8475 1.6050 0.9075 ;
        RECT 1.4400 0.4725 1.5000 0.5325 ;
        RECT 1.3350 0.8175 1.3950 0.8775 ;
        RECT 1.2225 0.4650 1.2825 0.5250 ;
        RECT 1.1250 0.1800 1.1850 0.2400 ;
        RECT 1.1250 0.8325 1.1850 0.8925 ;
        RECT 0.9150 0.1575 0.9750 0.2175 ;
        RECT 0.9150 0.8175 0.9750 0.8775 ;
        RECT 0.8100 0.4650 0.8700 0.5250 ;
        RECT 0.7050 0.6600 0.7650 0.7200 ;
        RECT 0.6000 0.4650 0.6600 0.5250 ;
        RECT 0.4950 0.1800 0.5550 0.2400 ;
        RECT 0.4950 0.8325 0.5550 0.8925 ;
        RECT 0.3825 0.4650 0.4425 0.5250 ;
        RECT 0.2850 0.6675 0.3450 0.7275 ;
        RECT 0.1725 0.4650 0.2325 0.5250 ;
        RECT 0.0750 0.1725 0.1350 0.2325 ;
        RECT 0.0750 0.8175 0.1350 0.8775 ;
        LAYER M1 ;
        RECT 1.6725 0.4650 1.9125 0.5850 ;
        RECT 1.5975 0.2625 1.6725 0.5850 ;
        RECT 1.4400 0.2625 1.5975 0.3375 ;
        RECT 1.4100 0.4125 1.5225 0.6975 ;
        RECT 1.3650 0.1500 1.4400 0.3375 ;
        RECT 1.3350 0.7950 1.4175 0.9000 ;
        RECT 1.3575 0.4125 1.4100 0.5700 ;
        RECT 1.0950 0.1500 1.3650 0.2550 ;
        RECT 1.2600 0.6450 1.3350 0.9000 ;
        RECT 1.0650 0.3450 1.2825 0.5700 ;
        RECT 0.8100 0.6450 1.2600 0.7200 ;
        RECT 0.8925 0.7950 0.9975 0.9000 ;
        RECT 0.8100 0.3375 0.9900 0.5550 ;
        RECT 0.1575 0.8250 0.8925 0.9000 ;
        RECT 0.4650 0.1575 0.8175 0.2625 ;
        RECT 0.7050 0.6300 0.8100 0.7500 ;
        RECT 0.5175 0.3375 0.7275 0.5550 ;
        RECT 0.2175 0.6450 0.6300 0.7500 ;
        RECT 0.3825 0.3375 0.4425 0.5700 ;
        RECT 0.3075 0.2100 0.3825 0.5700 ;
        RECT 0.0525 0.7950 0.1575 0.9000 ;
        LAYER VIA1 ;
        RECT 1.3650 0.1950 1.4400 0.2700 ;
        RECT 0.6975 0.1725 0.7725 0.2475 ;
        RECT 0.5175 0.6600 0.5925 0.7350 ;
        LAYER M2 ;
        RECT 1.3500 0.1125 1.4550 0.3075 ;
        RECT 0.7875 0.1125 1.3500 0.1875 ;
        RECT 0.7125 0.1125 0.7875 0.6975 ;
        RECT 0.6900 0.1125 0.7125 0.3000 ;
        RECT 0.6075 0.6225 0.7125 0.6975 ;
        RECT 0.5025 0.6225 0.6075 0.7725 ;
    END
END AO222_0011


MACRO AO222_0111
    CLASS CORE ;
    FOREIGN AO222_0111 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.7800 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 3.0975 0.2400 3.4125 0.7500 ;
        VIA 3.2550 0.3225 VIA12_slot ;
        VIA 3.2550 0.6675 VIA12_slot ;
        END
    END Z
    PIN C2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 2.1300 0.7125 2.5950 0.7875 ;
        RECT 2.0550 0.3600 2.1300 0.7875 ;
        VIA 2.0925 0.4725 VIA12_square ;
        END
    END C2
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 2.3625 0.5625 2.8275 0.6375 ;
        RECT 2.2875 0.4275 2.3625 0.6375 ;
        VIA 2.3250 0.5250 VIA12_square ;
        END
    END C1
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.6425 0.3600 1.7175 0.7875 ;
        RECT 1.1775 0.7125 1.6425 0.7875 ;
        VIA 1.6800 0.4500 VIA12_square ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.4100 0.4275 1.4850 0.6375 ;
        RECT 0.9450 0.5625 1.4100 0.6375 ;
        VIA 1.4475 0.5250 VIA12_square ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.8025 0.3300 0.8775 0.5700 ;
        RECT 0.2400 0.3300 0.8025 0.4050 ;
        RECT 0.1425 0.3300 0.2400 0.5550 ;
        RECT 0.0675 0.3300 0.1425 0.6825 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.5400 0.4050 0.6150 0.7875 ;
        RECT 0.0750 0.7125 0.5400 0.7875 ;
        VIA 0.5775 0.5250 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 3.7125 -0.0750 3.7800 0.0750 ;
        RECT 3.6375 -0.0750 3.7125 0.3150 ;
        RECT 3.3150 -0.0750 3.6375 0.0750 ;
        RECT 3.1950 -0.0750 3.3150 0.1950 ;
        RECT 2.8950 -0.0750 3.1950 0.0750 ;
        RECT 2.7750 -0.0750 2.8950 0.1950 ;
        RECT 2.0550 -0.0750 2.7750 0.0750 ;
        RECT 1.9350 -0.0750 2.0550 0.2475 ;
        RECT 1.8450 -0.0750 1.9350 0.0750 ;
        RECT 1.7250 -0.0750 1.8450 0.2475 ;
        RECT 1.0200 -0.0750 1.7250 0.0750 ;
        RECT 0.9150 -0.0750 1.0200 0.2550 ;
        RECT 0.1575 -0.0750 0.9150 0.0750 ;
        RECT 0.0525 -0.0750 0.1575 0.2475 ;
        RECT 0.0000 -0.0750 0.0525 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 3.7125 0.9750 3.7800 1.1250 ;
        RECT 3.6375 0.6375 3.7125 1.1250 ;
        RECT 3.3075 0.9750 3.6375 1.1250 ;
        RECT 3.2025 0.8025 3.3075 1.1250 ;
        RECT 2.8725 0.9750 3.2025 1.1250 ;
        RECT 2.7975 0.6375 2.8725 1.1250 ;
        RECT 2.4750 0.9750 2.7975 1.1250 ;
        RECT 2.3550 0.8025 2.4750 1.1250 ;
        RECT 2.0550 0.9750 2.3550 1.1250 ;
        RECT 1.9500 0.8025 2.0550 1.1250 ;
        RECT 0.0000 0.9750 1.9500 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 3.6450 0.2250 3.7050 0.2850 ;
        RECT 3.6450 0.6675 3.7050 0.7275 ;
        RECT 3.6450 0.8325 3.7050 0.8925 ;
        RECT 3.5400 0.4650 3.6000 0.5250 ;
        RECT 3.4350 0.2250 3.4950 0.2850 ;
        RECT 3.4350 0.7575 3.4950 0.8175 ;
        RECT 3.3300 0.4650 3.3900 0.5250 ;
        RECT 3.2250 0.1275 3.2850 0.1875 ;
        RECT 3.2250 0.8325 3.2850 0.8925 ;
        RECT 3.1200 0.4650 3.1800 0.5250 ;
        RECT 3.0150 0.2250 3.0750 0.2850 ;
        RECT 3.0150 0.7575 3.0750 0.8175 ;
        RECT 2.9100 0.4650 2.9700 0.5250 ;
        RECT 2.8050 0.1200 2.8650 0.1800 ;
        RECT 2.8050 0.6675 2.8650 0.7275 ;
        RECT 2.8050 0.8325 2.8650 0.8925 ;
        RECT 2.7000 0.4650 2.7600 0.5250 ;
        RECT 2.5950 0.6675 2.6550 0.7275 ;
        RECT 2.4900 0.4950 2.5500 0.5550 ;
        RECT 2.3850 0.1725 2.4450 0.2325 ;
        RECT 2.3850 0.8325 2.4450 0.8925 ;
        RECT 2.2800 0.4875 2.3400 0.5475 ;
        RECT 2.1750 0.6600 2.2350 0.7200 ;
        RECT 2.0700 0.4650 2.1300 0.5250 ;
        RECT 1.9650 0.1725 2.0250 0.2325 ;
        RECT 1.9650 0.8325 2.0250 0.8925 ;
        RECT 1.7550 0.1725 1.8150 0.2325 ;
        RECT 1.7550 0.8325 1.8150 0.8925 ;
        RECT 1.6500 0.4650 1.7100 0.5250 ;
        RECT 1.5450 0.6600 1.6050 0.7200 ;
        RECT 1.4400 0.4875 1.5000 0.5475 ;
        RECT 1.3350 0.1800 1.3950 0.2400 ;
        RECT 1.3350 0.8325 1.3950 0.8925 ;
        RECT 1.2300 0.4875 1.2900 0.5475 ;
        RECT 1.1250 0.6600 1.1850 0.7200 ;
        RECT 1.0200 0.4650 1.0800 0.5250 ;
        RECT 0.9150 0.1650 0.9750 0.2250 ;
        RECT 0.9150 0.8325 0.9750 0.8925 ;
        RECT 0.8100 0.4800 0.8700 0.5400 ;
        RECT 0.7050 0.6750 0.7650 0.7350 ;
        RECT 0.6000 0.4950 0.6600 0.5550 ;
        RECT 0.4950 0.1725 0.5550 0.2325 ;
        RECT 0.4950 0.8325 0.5550 0.8925 ;
        RECT 0.3900 0.4950 0.4500 0.5550 ;
        RECT 0.2850 0.6750 0.3450 0.7350 ;
        RECT 0.1800 0.4650 0.2400 0.5250 ;
        RECT 0.0750 0.1575 0.1350 0.2175 ;
        RECT 0.0750 0.8175 0.1350 0.8775 ;
        LAYER M1 ;
        RECT 2.9100 0.4425 3.6300 0.5475 ;
        RECT 3.4125 0.1950 3.5175 0.3675 ;
        RECT 3.4275 0.6225 3.5025 0.8700 ;
        RECT 3.0825 0.6225 3.4275 0.7125 ;
        RECT 3.0975 0.2775 3.4125 0.3675 ;
        RECT 2.9925 0.1950 3.0975 0.3675 ;
        RECT 3.0075 0.6225 3.0825 0.8700 ;
        RECT 2.8350 0.3000 2.9100 0.5475 ;
        RECT 2.6550 0.3225 2.7600 0.5550 ;
        RECT 1.0725 0.6525 2.6850 0.7275 ;
        RECT 2.1300 0.3225 2.6550 0.3975 ;
        RECT 2.2425 0.1500 2.5875 0.2475 ;
        RECT 2.2425 0.4725 2.5725 0.5775 ;
        RECT 2.0550 0.3225 2.1300 0.5550 ;
        RECT 0.1575 0.8250 1.8450 0.9000 ;
        RECT 1.6425 0.3300 1.7175 0.5550 ;
        RECT 1.0875 0.3300 1.6425 0.4050 ;
        RECT 1.2000 0.4800 1.5300 0.5775 ;
        RECT 1.2075 0.1500 1.5075 0.2550 ;
        RECT 1.0125 0.3300 1.0875 0.5625 ;
        RECT 0.4650 0.1500 0.8400 0.2550 ;
        RECT 0.2475 0.6600 0.8175 0.7425 ;
        RECT 0.3600 0.4800 0.6900 0.5775 ;
        RECT 0.0525 0.7950 0.1575 0.9000 ;
        LAYER VIA1 ;
        RECT 2.8350 0.3525 2.9100 0.4275 ;
        RECT 2.3775 0.1575 2.4525 0.2325 ;
        RECT 1.3275 0.1575 1.4025 0.2325 ;
        RECT 0.7050 0.1650 0.7800 0.2400 ;
        RECT 0.6975 0.6600 0.7725 0.7350 ;
        LAYER M2 ;
        RECT 2.8200 0.1575 2.9250 0.4650 ;
        RECT 1.3575 0.1575 2.8200 0.2325 ;
        RECT 1.2825 0.1125 1.3575 0.2325 ;
        RECT 0.7950 0.1125 1.2825 0.1875 ;
        RECT 0.6900 0.1125 0.7950 0.7800 ;
    END
END AO222_0111


MACRO AO222_1000
    CLASS CORE ;
    FOREIGN AO222_1000 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.8900 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 1.7775 0.1500 1.8525 0.9000 ;
        RECT 1.7475 0.1500 1.7775 0.3825 ;
        RECT 1.7325 0.6675 1.7775 0.9000 ;
        END
    END Z
    PIN C2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.2000 0.5625 1.6650 0.6375 ;
        VIA 1.4625 0.6000 VIA12_square ;
        END
    END C2
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.0575 0.4125 1.5225 0.4875 ;
        VIA 1.1700 0.4500 VIA12_square ;
        END
    END C1
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.9375 0.7125 1.4025 0.7875 ;
        RECT 0.8625 0.4050 0.9375 0.7875 ;
        VIA 0.9000 0.4875 VIA12_square ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.6150 0.3600 0.6375 0.5100 ;
        RECT 0.5325 0.1125 0.6150 0.5100 ;
        RECT 0.0675 0.1125 0.5325 0.1875 ;
        VIA 0.5850 0.4350 VIA12_square ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1425 0.4350 0.2325 0.5550 ;
        RECT 0.0675 0.3675 0.1425 0.6825 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.4275 0.8625 0.8925 0.9375 ;
        RECT 0.3525 0.4050 0.4275 0.9375 ;
        VIA 0.3900 0.4875 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.6350 -0.0750 1.8900 0.0750 ;
        RECT 1.5150 -0.0750 1.6350 0.1800 ;
        RECT 0.9975 -0.0750 1.5150 0.0750 ;
        RECT 0.8925 -0.0750 0.9975 0.2400 ;
        RECT 0.1425 -0.0750 0.8925 0.0750 ;
        RECT 0.0675 -0.0750 0.1425 0.2625 ;
        RECT 0.0000 -0.0750 0.0675 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.6350 0.9750 1.8900 1.1250 ;
        RECT 1.5150 0.8250 1.6350 1.1250 ;
        RECT 1.1850 0.9750 1.5150 1.1250 ;
        RECT 1.0800 0.8025 1.1850 1.1250 ;
        RECT 0.0000 0.9750 1.0800 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.7550 0.1800 1.8150 0.2400 ;
        RECT 1.7550 0.8175 1.8150 0.8775 ;
        RECT 1.6425 0.4950 1.7025 0.5550 ;
        RECT 1.5450 0.1200 1.6050 0.1800 ;
        RECT 1.5450 0.8475 1.6050 0.9075 ;
        RECT 1.4400 0.4725 1.5000 0.5325 ;
        RECT 1.3350 0.8175 1.3950 0.8775 ;
        RECT 1.2225 0.4650 1.2825 0.5250 ;
        RECT 1.1250 0.1800 1.1850 0.2400 ;
        RECT 1.1250 0.8325 1.1850 0.8925 ;
        RECT 0.9150 0.1575 0.9750 0.2175 ;
        RECT 0.9150 0.8175 0.9750 0.8775 ;
        RECT 0.8100 0.4650 0.8700 0.5250 ;
        RECT 0.7050 0.6600 0.7650 0.7200 ;
        RECT 0.6000 0.4650 0.6600 0.5250 ;
        RECT 0.4950 0.1800 0.5550 0.2400 ;
        RECT 0.4950 0.8325 0.5550 0.8925 ;
        RECT 0.3825 0.4650 0.4425 0.5250 ;
        RECT 0.2850 0.6675 0.3450 0.7275 ;
        RECT 0.1725 0.4650 0.2325 0.5250 ;
        RECT 0.0750 0.1575 0.1350 0.2175 ;
        RECT 0.0750 0.8175 0.1350 0.8775 ;
        LAYER M1 ;
        RECT 1.6725 0.4650 1.7025 0.5850 ;
        RECT 1.5975 0.2625 1.6725 0.5850 ;
        RECT 1.4400 0.2625 1.5975 0.3375 ;
        RECT 1.4100 0.4125 1.5225 0.6975 ;
        RECT 1.3650 0.1500 1.4400 0.3375 ;
        RECT 1.3350 0.7950 1.4175 0.9000 ;
        RECT 1.3575 0.4125 1.4100 0.5700 ;
        RECT 1.0950 0.1500 1.3650 0.2550 ;
        RECT 1.2600 0.6450 1.3350 0.9000 ;
        RECT 1.0650 0.3450 1.2825 0.5700 ;
        RECT 0.8100 0.6450 1.2600 0.7200 ;
        RECT 0.8925 0.7950 0.9975 0.9000 ;
        RECT 0.8100 0.3375 0.9900 0.5550 ;
        RECT 0.1575 0.8250 0.8925 0.9000 ;
        RECT 0.4650 0.1575 0.8175 0.2625 ;
        RECT 0.7050 0.6300 0.8100 0.7500 ;
        RECT 0.5175 0.3375 0.7275 0.5550 ;
        RECT 0.2175 0.6450 0.6300 0.7500 ;
        RECT 0.3825 0.3375 0.4425 0.5700 ;
        RECT 0.3075 0.2100 0.3825 0.5700 ;
        RECT 0.0525 0.7950 0.1575 0.9000 ;
        LAYER VIA1 ;
        RECT 1.3650 0.1950 1.4400 0.2700 ;
        RECT 0.6975 0.1725 0.7725 0.2475 ;
        RECT 0.5175 0.6600 0.5925 0.7350 ;
        LAYER M2 ;
        RECT 1.3500 0.1125 1.4550 0.3075 ;
        RECT 0.7875 0.1125 1.3500 0.1875 ;
        RECT 0.7125 0.1125 0.7875 0.6975 ;
        RECT 0.6900 0.1125 0.7125 0.3000 ;
        RECT 0.6075 0.6225 0.7125 0.6975 ;
        RECT 0.5025 0.6225 0.6075 0.7725 ;
    END
END AO222_1000


MACRO AO222_1010
    CLASS CORE ;
    FOREIGN AO222_1010 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.8900 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 1.7775 0.2175 1.8525 0.8325 ;
        RECT 1.7475 0.2175 1.7775 0.3825 ;
        RECT 1.7475 0.6675 1.7775 0.8325 ;
        END
    END Z
    PIN C2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.2000 0.5625 1.6650 0.6375 ;
        VIA 1.4625 0.6000 VIA12_square ;
        END
    END C2
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.0575 0.4125 1.5225 0.4875 ;
        VIA 1.1700 0.4500 VIA12_square ;
        END
    END C1
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.9375 0.7125 1.4025 0.7875 ;
        RECT 0.8625 0.4050 0.9375 0.7875 ;
        VIA 0.9000 0.4875 VIA12_square ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.6150 0.3600 0.6375 0.5100 ;
        RECT 0.5325 0.1125 0.6150 0.5100 ;
        RECT 0.0675 0.1125 0.5325 0.1875 ;
        VIA 0.5850 0.4350 VIA12_square ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1425 0.4350 0.2325 0.5550 ;
        RECT 0.0675 0.3675 0.1425 0.6825 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.4275 0.8625 0.8925 0.9375 ;
        RECT 0.3525 0.4050 0.4275 0.9375 ;
        VIA 0.3900 0.4875 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.6350 -0.0750 1.8900 0.0750 ;
        RECT 1.5150 -0.0750 1.6350 0.1800 ;
        RECT 0.9975 -0.0750 1.5150 0.0750 ;
        RECT 0.8925 -0.0750 0.9975 0.2400 ;
        RECT 0.1425 -0.0750 0.8925 0.0750 ;
        RECT 0.0675 -0.0750 0.1425 0.2625 ;
        RECT 0.0000 -0.0750 0.0675 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.6350 0.9750 1.8900 1.1250 ;
        RECT 1.5150 0.8250 1.6350 1.1250 ;
        RECT 1.1850 0.9750 1.5150 1.1250 ;
        RECT 1.0800 0.8025 1.1850 1.1250 ;
        RECT 0.0000 0.9750 1.0800 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.7550 0.2700 1.8150 0.3300 ;
        RECT 1.7550 0.7200 1.8150 0.7800 ;
        RECT 1.6425 0.4950 1.7025 0.5550 ;
        RECT 1.5450 0.1200 1.6050 0.1800 ;
        RECT 1.5450 0.8475 1.6050 0.9075 ;
        RECT 1.4400 0.4725 1.5000 0.5325 ;
        RECT 1.3350 0.8175 1.3950 0.8775 ;
        RECT 1.2225 0.4650 1.2825 0.5250 ;
        RECT 1.1250 0.1800 1.1850 0.2400 ;
        RECT 1.1250 0.8325 1.1850 0.8925 ;
        RECT 0.9150 0.1575 0.9750 0.2175 ;
        RECT 0.9150 0.8175 0.9750 0.8775 ;
        RECT 0.8100 0.4650 0.8700 0.5250 ;
        RECT 0.7050 0.6600 0.7650 0.7200 ;
        RECT 0.6000 0.4650 0.6600 0.5250 ;
        RECT 0.4950 0.1800 0.5550 0.2400 ;
        RECT 0.4950 0.8325 0.5550 0.8925 ;
        RECT 0.3825 0.4650 0.4425 0.5250 ;
        RECT 0.2850 0.6675 0.3450 0.7275 ;
        RECT 0.1725 0.4650 0.2325 0.5250 ;
        RECT 0.0750 0.1725 0.1350 0.2325 ;
        RECT 0.0750 0.8175 0.1350 0.8775 ;
        LAYER M1 ;
        RECT 1.6725 0.4650 1.7025 0.5850 ;
        RECT 1.5975 0.2625 1.6725 0.5850 ;
        RECT 1.4400 0.2625 1.5975 0.3375 ;
        RECT 1.4100 0.4125 1.5225 0.6975 ;
        RECT 1.3650 0.1500 1.4400 0.3375 ;
        RECT 1.3350 0.7950 1.4175 0.9000 ;
        RECT 1.3575 0.4125 1.4100 0.5700 ;
        RECT 1.0950 0.1500 1.3650 0.2550 ;
        RECT 1.2600 0.6450 1.3350 0.9000 ;
        RECT 1.0650 0.3450 1.2825 0.5700 ;
        RECT 0.8100 0.6450 1.2600 0.7200 ;
        RECT 0.8925 0.7950 0.9975 0.9000 ;
        RECT 0.8100 0.3375 0.9900 0.5550 ;
        RECT 0.1575 0.8250 0.8925 0.9000 ;
        RECT 0.4650 0.1575 0.8175 0.2625 ;
        RECT 0.7050 0.6300 0.8100 0.7500 ;
        RECT 0.5175 0.3375 0.7275 0.5550 ;
        RECT 0.2175 0.6450 0.6300 0.7500 ;
        RECT 0.3825 0.3375 0.4425 0.5700 ;
        RECT 0.3075 0.2100 0.3825 0.5700 ;
        RECT 0.0525 0.7950 0.1575 0.9000 ;
        LAYER VIA1 ;
        RECT 1.3650 0.1950 1.4400 0.2700 ;
        RECT 0.6975 0.1725 0.7725 0.2475 ;
        RECT 0.5175 0.6600 0.5925 0.7350 ;
        LAYER M2 ;
        RECT 1.3500 0.1125 1.4550 0.3075 ;
        RECT 0.7875 0.1125 1.3500 0.1875 ;
        RECT 0.7125 0.1125 0.7875 0.6975 ;
        RECT 0.6900 0.1125 0.7125 0.3000 ;
        RECT 0.6075 0.6225 0.7125 0.6975 ;
        RECT 0.5025 0.6225 0.6075 0.7725 ;
    END
END AO222_1010


MACRO AO22_0011
    CLASS CORE ;
    FOREIGN AO22_0011 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.6800 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 1.5675 0.3075 1.6425 0.7425 ;
        RECT 1.4025 0.3075 1.5675 0.3825 ;
        RECT 1.4025 0.6675 1.5675 0.7425 ;
        RECT 1.3275 0.2175 1.4025 0.3825 ;
        RECT 1.3275 0.6675 1.4025 0.8550 ;
        END
    END Z
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.8625 0.5625 1.3275 0.6375 ;
        VIA 0.9750 0.6000 VIA12_square ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.7425 0.8625 1.2075 0.9375 ;
        RECT 0.6375 0.5400 0.7425 0.9375 ;
        RECT 0.5925 0.5400 0.6375 0.6450 ;
        VIA 0.6675 0.5925 VIA12_square ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1425 0.4050 0.2700 0.5100 ;
        RECT 0.0675 0.3675 0.1425 0.6825 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.6075 0.2625 1.0950 0.3375 ;
        RECT 0.5025 0.2625 0.6075 0.4350 ;
        VIA 0.5475 0.3525 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.6350 -0.0750 1.6800 0.0750 ;
        RECT 1.5150 -0.0750 1.6350 0.2175 ;
        RECT 1.2150 -0.0750 1.5150 0.0750 ;
        RECT 1.0950 -0.0750 1.2150 0.2175 ;
        RECT 1.0050 -0.0750 1.0950 0.0750 ;
        RECT 0.8850 -0.0750 1.0050 0.2175 ;
        RECT 0.1575 -0.0750 0.8850 0.0750 ;
        RECT 0.0450 -0.0750 0.1575 0.2475 ;
        RECT 0.0000 -0.0750 0.0450 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.6350 0.9750 1.6800 1.1250 ;
        RECT 1.5150 0.8175 1.6350 1.1250 ;
        RECT 1.2150 0.9750 1.5150 1.1250 ;
        RECT 1.0950 0.8025 1.2150 1.1250 ;
        RECT 0.7950 0.9750 1.0950 1.1250 ;
        RECT 0.6750 0.8700 0.7950 1.1250 ;
        RECT 0.0000 0.9750 0.6750 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.5450 0.1575 1.6050 0.2175 ;
        RECT 1.5450 0.8325 1.6050 0.8925 ;
        RECT 1.4325 0.4950 1.4925 0.5550 ;
        RECT 1.3350 0.2700 1.3950 0.3300 ;
        RECT 1.3350 0.7650 1.3950 0.8250 ;
        RECT 1.2300 0.4950 1.2900 0.5550 ;
        RECT 1.1250 0.1575 1.1850 0.2175 ;
        RECT 1.1250 0.8325 1.1850 0.8925 ;
        RECT 0.9150 0.1575 0.9750 0.2175 ;
        RECT 0.9150 0.7575 0.9750 0.8175 ;
        RECT 0.8175 0.4950 0.8775 0.5550 ;
        RECT 0.7050 0.8700 0.7650 0.9300 ;
        RECT 0.6000 0.4950 0.6600 0.5550 ;
        RECT 0.4950 0.1575 0.5550 0.2175 ;
        RECT 0.4950 0.8325 0.5550 0.8925 ;
        RECT 0.3825 0.4500 0.4425 0.5100 ;
        RECT 0.2850 0.6525 0.3450 0.7125 ;
        RECT 0.0750 0.1575 0.1350 0.2175 ;
        RECT 0.0750 0.8250 0.1350 0.8850 ;
        RECT 0.1800 0.4500 0.2400 0.5100 ;
        LAYER M1 ;
        RECT 1.2525 0.4650 1.4925 0.5850 ;
        RECT 1.1775 0.2925 1.2525 0.5850 ;
        RECT 0.8100 0.2925 1.1775 0.3675 ;
        RECT 0.8175 0.4500 1.0875 0.6375 ;
        RECT 0.8850 0.7200 0.9750 0.8550 ;
        RECT 0.6000 0.7200 0.8850 0.7950 ;
        RECT 0.7350 0.1500 0.8100 0.3675 ;
        RECT 0.5475 0.4800 0.7425 0.6450 ;
        RECT 0.2625 0.1500 0.7350 0.2325 ;
        RECT 0.4725 0.3075 0.6300 0.4050 ;
        RECT 0.5250 0.7200 0.6000 0.9000 ;
        RECT 0.1500 0.8250 0.5250 0.9000 ;
        RECT 0.3525 0.3075 0.4725 0.5100 ;
        RECT 0.2175 0.5850 0.4500 0.7500 ;
        RECT 0.0450 0.7950 0.1500 0.9000 ;
        LAYER VIA1 ;
        RECT 0.3525 0.6300 0.4275 0.7050 ;
        RECT 0.3075 0.1575 0.3825 0.2325 ;
        LAYER M2 ;
        RECT 0.3525 0.1575 0.4275 0.7500 ;
        RECT 0.2625 0.1575 0.3525 0.2325 ;
    END
END AO22_0011


MACRO AO22_0111
    CLASS CORE ;
    FOREIGN AO22_0111 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.9400 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 2.2575 0.2400 2.5725 0.7500 ;
        VIA 2.4150 0.3225 VIA12_slot ;
        VIA 2.4150 0.6675 VIA12_slot ;
        END
    END Z
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.2900 0.7125 1.7550 0.7875 ;
        RECT 1.2150 0.3600 1.2900 0.7875 ;
        VIA 1.2525 0.4725 VIA12_square ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.5225 0.5625 1.9875 0.6375 ;
        RECT 1.4475 0.4275 1.5225 0.6375 ;
        VIA 1.4850 0.5250 VIA12_square ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.8025 0.3300 0.8775 0.5700 ;
        RECT 0.2400 0.3300 0.8025 0.4050 ;
        RECT 0.1425 0.3300 0.2400 0.5550 ;
        RECT 0.0675 0.3300 0.1425 0.6825 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.5400 0.4050 0.6150 0.7875 ;
        RECT 0.0750 0.7125 0.5400 0.7875 ;
        VIA 0.5775 0.5250 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 2.8725 -0.0750 2.9400 0.0750 ;
        RECT 2.7975 -0.0750 2.8725 0.3150 ;
        RECT 2.4750 -0.0750 2.7975 0.0750 ;
        RECT 2.3550 -0.0750 2.4750 0.1950 ;
        RECT 2.0550 -0.0750 2.3550 0.0750 ;
        RECT 1.9350 -0.0750 2.0550 0.1950 ;
        RECT 1.2150 -0.0750 1.9350 0.0750 ;
        RECT 1.0950 -0.0750 1.2150 0.2475 ;
        RECT 1.0200 -0.0750 1.0950 0.0750 ;
        RECT 0.9150 -0.0750 1.0200 0.2550 ;
        RECT 0.1575 -0.0750 0.9150 0.0750 ;
        RECT 0.0525 -0.0750 0.1575 0.2475 ;
        RECT 0.0000 -0.0750 0.0525 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 2.8725 0.9750 2.9400 1.1250 ;
        RECT 2.7975 0.6375 2.8725 1.1250 ;
        RECT 2.4675 0.9750 2.7975 1.1250 ;
        RECT 2.3625 0.8025 2.4675 1.1250 ;
        RECT 2.0325 0.9750 2.3625 1.1250 ;
        RECT 1.9575 0.6375 2.0325 1.1250 ;
        RECT 1.6350 0.9750 1.9575 1.1250 ;
        RECT 1.5150 0.8025 1.6350 1.1250 ;
        RECT 1.2150 0.9750 1.5150 1.1250 ;
        RECT 1.1100 0.8025 1.2150 1.1250 ;
        RECT 0.0000 0.9750 1.1100 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 2.8050 0.2250 2.8650 0.2850 ;
        RECT 2.8050 0.6675 2.8650 0.7275 ;
        RECT 2.8050 0.8325 2.8650 0.8925 ;
        RECT 2.7000 0.4650 2.7600 0.5250 ;
        RECT 2.5950 0.2250 2.6550 0.2850 ;
        RECT 2.5950 0.7575 2.6550 0.8175 ;
        RECT 2.4900 0.4650 2.5500 0.5250 ;
        RECT 2.3850 0.1275 2.4450 0.1875 ;
        RECT 2.3850 0.8325 2.4450 0.8925 ;
        RECT 2.2800 0.4650 2.3400 0.5250 ;
        RECT 2.1750 0.2250 2.2350 0.2850 ;
        RECT 2.1750 0.7575 2.2350 0.8175 ;
        RECT 2.0700 0.4650 2.1300 0.5250 ;
        RECT 1.9650 0.1200 2.0250 0.1800 ;
        RECT 1.9650 0.6675 2.0250 0.7275 ;
        RECT 1.9650 0.8325 2.0250 0.8925 ;
        RECT 1.8600 0.4650 1.9200 0.5250 ;
        RECT 1.7550 0.6675 1.8150 0.7275 ;
        RECT 1.6500 0.4950 1.7100 0.5550 ;
        RECT 1.5450 0.1725 1.6050 0.2325 ;
        RECT 1.5450 0.8325 1.6050 0.8925 ;
        RECT 1.4400 0.4875 1.5000 0.5475 ;
        RECT 1.3350 0.6600 1.3950 0.7200 ;
        RECT 1.2300 0.4650 1.2900 0.5250 ;
        RECT 1.1250 0.1725 1.1850 0.2325 ;
        RECT 1.1250 0.8325 1.1850 0.8925 ;
        RECT 0.9150 0.1650 0.9750 0.2250 ;
        RECT 0.9150 0.8325 0.9750 0.8925 ;
        RECT 0.8100 0.4800 0.8700 0.5400 ;
        RECT 0.7050 0.6750 0.7650 0.7350 ;
        RECT 0.6000 0.4950 0.6600 0.5550 ;
        RECT 0.4950 0.1725 0.5550 0.2325 ;
        RECT 0.4950 0.8325 0.5550 0.8925 ;
        RECT 0.3900 0.4950 0.4500 0.5550 ;
        RECT 0.2850 0.6750 0.3450 0.7350 ;
        RECT 0.1800 0.4650 0.2400 0.5250 ;
        RECT 0.0750 0.1575 0.1350 0.2175 ;
        RECT 0.0750 0.8175 0.1350 0.8775 ;
        LAYER M1 ;
        RECT 2.0700 0.4425 2.7900 0.5475 ;
        RECT 2.5725 0.1950 2.6775 0.3675 ;
        RECT 2.5875 0.6225 2.6625 0.8700 ;
        RECT 2.2425 0.6225 2.5875 0.7125 ;
        RECT 2.2575 0.2775 2.5725 0.3675 ;
        RECT 2.1525 0.1950 2.2575 0.3675 ;
        RECT 2.1675 0.6225 2.2425 0.8700 ;
        RECT 1.9950 0.3000 2.0700 0.5475 ;
        RECT 1.8150 0.3225 1.9200 0.5550 ;
        RECT 1.0050 0.6525 1.8450 0.7275 ;
        RECT 1.2900 0.3225 1.8150 0.3975 ;
        RECT 1.4025 0.1500 1.7475 0.2475 ;
        RECT 1.4025 0.4725 1.7325 0.5775 ;
        RECT 1.2150 0.3225 1.2900 0.5550 ;
        RECT 0.9225 0.6525 1.0050 0.9000 ;
        RECT 0.1575 0.8250 0.9225 0.9000 ;
        RECT 0.4650 0.1500 0.8400 0.2550 ;
        RECT 0.2475 0.6600 0.8175 0.7425 ;
        RECT 0.3600 0.4800 0.6900 0.5775 ;
        RECT 0.0525 0.7950 0.1575 0.9000 ;
        LAYER VIA1 ;
        RECT 1.9950 0.3525 2.0700 0.4275 ;
        RECT 1.5375 0.1575 1.6125 0.2325 ;
        RECT 0.7050 0.1650 0.7800 0.2400 ;
        RECT 0.6975 0.6600 0.7725 0.7350 ;
        LAYER M2 ;
        RECT 1.9800 0.1575 2.0850 0.4650 ;
        RECT 1.5675 0.1575 1.9800 0.2325 ;
        RECT 1.4925 0.1125 1.5675 0.2325 ;
        RECT 0.7950 0.1125 1.4925 0.1875 ;
        RECT 0.6900 0.1125 0.7950 0.7800 ;
    END
END AO22_0111


MACRO AO22_1000
    CLASS CORE ;
    FOREIGN AO22_1000 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.4700 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 1.3575 0.1500 1.4325 0.9000 ;
        RECT 1.3275 0.1500 1.3575 0.3825 ;
        RECT 1.3125 0.6675 1.3575 0.9000 ;
        END
    END Z
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.8625 0.5625 1.3275 0.6375 ;
        VIA 0.9750 0.6000 VIA12_square ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.7425 0.8625 1.2075 0.9375 ;
        RECT 0.6375 0.5400 0.7425 0.9375 ;
        RECT 0.5925 0.5400 0.6375 0.6450 ;
        VIA 0.6675 0.5925 VIA12_square ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1425 0.4050 0.2700 0.5100 ;
        RECT 0.0675 0.3675 0.1425 0.6825 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.6075 0.2625 1.0950 0.3375 ;
        RECT 0.5025 0.2625 0.6075 0.4350 ;
        VIA 0.5475 0.3525 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.2150 -0.0750 1.4700 0.0750 ;
        RECT 1.0950 -0.0750 1.2150 0.2175 ;
        RECT 1.0050 -0.0750 1.0950 0.0750 ;
        RECT 0.8850 -0.0750 1.0050 0.2175 ;
        RECT 0.1575 -0.0750 0.8850 0.0750 ;
        RECT 0.0450 -0.0750 0.1575 0.2475 ;
        RECT 0.0000 -0.0750 0.0450 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.2150 0.9750 1.4700 1.1250 ;
        RECT 1.0950 0.8025 1.2150 1.1250 ;
        RECT 0.7950 0.9750 1.0950 1.1250 ;
        RECT 0.6750 0.8700 0.7950 1.1250 ;
        RECT 0.0000 0.9750 0.6750 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.3350 0.1800 1.3950 0.2400 ;
        RECT 1.3350 0.8175 1.3950 0.8775 ;
        RECT 1.2225 0.4725 1.2825 0.5325 ;
        RECT 1.1250 0.1575 1.1850 0.2175 ;
        RECT 1.1250 0.8325 1.1850 0.8925 ;
        RECT 0.9150 0.1575 0.9750 0.2175 ;
        RECT 0.9150 0.8175 0.9750 0.8775 ;
        RECT 0.8175 0.4950 0.8775 0.5550 ;
        RECT 0.7050 0.8700 0.7650 0.9300 ;
        RECT 0.6000 0.4950 0.6600 0.5550 ;
        RECT 0.4950 0.1575 0.5550 0.2175 ;
        RECT 0.3825 0.4500 0.4425 0.5100 ;
        RECT 0.2850 0.6525 0.3450 0.7125 ;
        RECT 0.1800 0.4500 0.2400 0.5100 ;
        RECT 0.0750 0.1575 0.1350 0.2175 ;
        RECT 0.0750 0.8250 0.1350 0.8850 ;
        RECT 0.4950 0.8325 0.5550 0.8925 ;
        LAYER M1 ;
        RECT 1.2525 0.4425 1.2825 0.5625 ;
        RECT 1.1775 0.2925 1.2525 0.5625 ;
        RECT 0.8100 0.2925 1.1775 0.3675 ;
        RECT 0.8175 0.4500 1.0875 0.6375 ;
        RECT 0.8850 0.7200 0.9975 0.9000 ;
        RECT 0.6000 0.7200 0.8850 0.7950 ;
        RECT 0.7350 0.1500 0.8100 0.3675 ;
        RECT 0.5475 0.4800 0.7425 0.6450 ;
        RECT 0.2625 0.1500 0.7350 0.2325 ;
        RECT 0.4725 0.3075 0.6300 0.4050 ;
        RECT 0.5250 0.7200 0.6000 0.9000 ;
        RECT 0.1500 0.8250 0.5250 0.9000 ;
        RECT 0.3525 0.3075 0.4725 0.5100 ;
        RECT 0.2175 0.5850 0.4500 0.7500 ;
        RECT 0.0450 0.7950 0.1500 0.9000 ;
        LAYER VIA1 ;
        RECT 0.3525 0.6300 0.4275 0.7050 ;
        RECT 0.3075 0.1575 0.3825 0.2325 ;
        LAYER M2 ;
        RECT 0.3525 0.1575 0.4275 0.7500 ;
        RECT 0.2625 0.1575 0.3525 0.2325 ;
    END
END AO22_1000


MACRO AO22_1010
    CLASS CORE ;
    FOREIGN AO22_1010 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.4700 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 1.3575 0.2175 1.4325 0.8325 ;
        RECT 1.3275 0.2175 1.3575 0.3825 ;
        RECT 1.3275 0.6675 1.3575 0.8325 ;
        END
    END Z
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.8925 0.5625 1.3575 0.6375 ;
        VIA 1.0050 0.6000 VIA12_square ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.6975 0.7125 1.1175 0.7875 ;
        RECT 0.5925 0.5100 0.6975 0.7875 ;
        VIA 0.6450 0.5925 VIA12_square ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1425 0.4050 0.2700 0.5100 ;
        RECT 0.0675 0.3675 0.1425 0.6825 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.6075 0.2625 0.9675 0.3375 ;
        RECT 0.5025 0.2625 0.6075 0.4350 ;
        VIA 0.5550 0.3525 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.2150 -0.0750 1.4700 0.0750 ;
        RECT 1.0950 -0.0750 1.2150 0.2175 ;
        RECT 1.0050 -0.0750 1.0950 0.0750 ;
        RECT 0.8850 -0.0750 1.0050 0.2175 ;
        RECT 0.1575 -0.0750 0.8850 0.0750 ;
        RECT 0.0450 -0.0750 0.1575 0.2475 ;
        RECT 0.0000 -0.0750 0.0450 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.2150 0.9750 1.4700 1.1250 ;
        RECT 1.0950 0.8025 1.2150 1.1250 ;
        RECT 0.7950 0.9750 1.0950 1.1250 ;
        RECT 0.6750 0.8700 0.7950 1.1250 ;
        RECT 0.0000 0.9750 0.6750 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.3350 0.2700 1.3950 0.3300 ;
        RECT 1.3350 0.7200 1.3950 0.7800 ;
        RECT 1.2225 0.4725 1.2825 0.5325 ;
        RECT 1.1250 0.1575 1.1850 0.2175 ;
        RECT 1.1250 0.8325 1.1850 0.8925 ;
        RECT 0.9150 0.1575 0.9750 0.2175 ;
        RECT 0.9150 0.7575 0.9750 0.8175 ;
        RECT 0.8175 0.4950 0.8775 0.5550 ;
        RECT 0.7050 0.8700 0.7650 0.9300 ;
        RECT 0.6000 0.4950 0.6600 0.5550 ;
        RECT 0.4950 0.1650 0.5550 0.2250 ;
        RECT 0.4950 0.8325 0.5550 0.8925 ;
        RECT 0.3825 0.4500 0.4425 0.5100 ;
        RECT 0.2850 0.6525 0.3450 0.7125 ;
        RECT 0.0750 0.1575 0.1350 0.2175 ;
        RECT 0.0750 0.8250 0.1350 0.8850 ;
        RECT 0.1800 0.4500 0.2400 0.5100 ;
        LAYER M1 ;
        RECT 1.2525 0.4425 1.2825 0.5625 ;
        RECT 1.1775 0.2925 1.2525 0.5625 ;
        RECT 0.8100 0.2925 1.1775 0.3675 ;
        RECT 0.8175 0.4500 1.0875 0.6375 ;
        RECT 0.8850 0.7200 0.9750 0.8550 ;
        RECT 0.6000 0.7200 0.8850 0.7950 ;
        RECT 0.7350 0.1500 0.8100 0.3675 ;
        RECT 0.5475 0.4800 0.7425 0.6450 ;
        RECT 0.4275 0.1500 0.7350 0.2250 ;
        RECT 0.4800 0.3000 0.6300 0.4050 ;
        RECT 0.5250 0.7200 0.6000 0.9000 ;
        RECT 0.1500 0.8250 0.5250 0.9000 ;
        RECT 0.4725 0.3075 0.4800 0.4050 ;
        RECT 0.3525 0.3075 0.4725 0.5100 ;
        RECT 0.2550 0.5850 0.4500 0.7500 ;
        RECT 0.2625 0.1500 0.4275 0.2325 ;
        RECT 0.0450 0.7950 0.1500 0.9000 ;
        LAYER VIA1 ;
        RECT 0.3675 0.6300 0.4425 0.7050 ;
        RECT 0.3075 0.1575 0.3825 0.2325 ;
        LAYER M2 ;
        RECT 0.4275 0.5850 0.4575 0.7425 ;
        RECT 0.3525 0.1575 0.4275 0.7425 ;
        RECT 0.2625 0.1575 0.3525 0.2325 ;
    END
END AO22_1010


MACRO AO31_0011
    CLASS CORE ;
    FOREIGN AO31_0011 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.4700 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 1.3575 0.3150 1.4325 0.7425 ;
        RECT 1.1925 0.3150 1.3575 0.3900 ;
        RECT 1.1925 0.6675 1.3575 0.7425 ;
        RECT 1.1175 0.2175 1.1925 0.3900 ;
        RECT 1.1175 0.6675 1.1925 0.8550 ;
        END
    END Z
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.8475 0.1125 1.1925 0.1875 ;
        RECT 0.7725 0.1125 0.8475 0.5250 ;
        RECT 0.6525 0.1125 0.7725 0.1875 ;
        VIA 0.8100 0.4425 VIA12_square ;
        END
    END B
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.0675 0.2625 0.5325 0.3375 ;
        VIA 0.2550 0.3000 VIA12_square ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.4725 0.8625 0.9225 0.9375 ;
        RECT 0.3675 0.4350 0.4725 0.9375 ;
        VIA 0.4200 0.5175 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.6525 0.7125 1.0875 0.7875 ;
        RECT 0.5775 0.3975 0.6525 0.7875 ;
        VIA 0.6150 0.5175 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.4250 -0.0750 1.4700 0.0750 ;
        RECT 1.3050 -0.0750 1.4250 0.2175 ;
        RECT 1.0050 -0.0750 1.3050 0.0750 ;
        RECT 0.8850 -0.0750 1.0050 0.1800 ;
        RECT 0.1425 -0.0750 0.8850 0.0750 ;
        RECT 0.0675 -0.0750 0.1425 0.3225 ;
        RECT 0.0000 -0.0750 0.0675 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.4250 0.9750 1.4700 1.1250 ;
        RECT 1.3050 0.8175 1.4250 1.1250 ;
        RECT 1.0050 0.9750 1.3050 1.1250 ;
        RECT 0.9000 0.8400 1.0050 1.1250 ;
        RECT 0.0000 0.9750 0.9000 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.3350 0.1575 1.3950 0.2175 ;
        RECT 1.3350 0.8325 1.3950 0.8925 ;
        RECT 1.2225 0.4950 1.2825 0.5550 ;
        RECT 1.1250 0.2550 1.1850 0.3150 ;
        RECT 1.1250 0.7650 1.1850 0.8250 ;
        RECT 1.0200 0.4950 1.0800 0.5550 ;
        RECT 0.9150 0.1200 0.9750 0.1800 ;
        RECT 0.9150 0.8700 0.9750 0.9300 ;
        RECT 0.8100 0.4800 0.8700 0.5400 ;
        RECT 0.7050 0.2400 0.7650 0.3000 ;
        RECT 0.7050 0.8325 0.7650 0.8925 ;
        RECT 0.5925 0.4950 0.6525 0.5550 ;
        RECT 0.4950 0.6825 0.5550 0.7425 ;
        RECT 0.3900 0.4875 0.4500 0.5475 ;
        RECT 0.2850 0.8325 0.3450 0.8925 ;
        RECT 0.1800 0.4950 0.2400 0.5550 ;
        RECT 0.0750 0.2250 0.1350 0.2850 ;
        RECT 0.0750 0.7575 0.1350 0.8175 ;
        LAYER M1 ;
        RECT 1.0425 0.4650 1.2825 0.5850 ;
        RECT 0.9675 0.2550 1.0425 0.7500 ;
        RECT 0.7725 0.2550 0.9675 0.3300 ;
        RECT 0.1425 0.6750 0.9675 0.7500 ;
        RECT 0.7275 0.4050 0.8925 0.6000 ;
        RECT 0.2550 0.8250 0.7950 0.9000 ;
        RECT 0.6975 0.2100 0.7725 0.3300 ;
        RECT 0.6225 0.4275 0.6525 0.6000 ;
        RECT 0.5475 0.2175 0.6225 0.6000 ;
        RECT 0.3675 0.2175 0.4725 0.6000 ;
        RECT 0.2175 0.2175 0.2925 0.5850 ;
        RECT 0.1725 0.4650 0.2175 0.5850 ;
        RECT 0.0675 0.6750 0.1425 0.8475 ;
    END
END AO31_0011


MACRO AO31_0111
    CLASS CORE ;
    FOREIGN AO31_0111 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.7300 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 1.8375 0.3000 2.1525 0.7725 ;
        VIA 1.9950 0.3600 VIA12_slot ;
        VIA 1.9950 0.7125 VIA12_slot ;
        END
    END Z
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 2.3775 0.4125 2.6325 0.4875 ;
        RECT 2.3025 0.1125 2.3775 0.4875 ;
        RECT 1.6425 0.1125 2.3025 0.1875 ;
        RECT 1.5675 0.1125 1.6425 0.4875 ;
        RECT 1.5225 0.4125 1.5675 0.4875 ;
        RECT 1.4175 0.4125 1.5225 0.6075 ;
        VIA 2.5500 0.4500 VIA12_square ;
        VIA 1.4700 0.5325 VIA12_square ;
        END
    END B
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.6825 0.5625 1.1100 0.6375 ;
        RECT 0.5775 0.4725 0.6825 0.6375 ;
        VIA 0.6300 0.5475 VIA12_square ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.8025 0.4125 1.2675 0.4875 ;
        VIA 1.0275 0.4500 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.1425 0.2625 1.3050 0.3375 ;
        VIA 1.1925 0.3000 VIA12_square ;
        VIA 0.2550 0.3000 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 2.4750 -0.0750 2.7300 0.0750 ;
        RECT 2.3550 -0.0750 2.4750 0.1800 ;
        RECT 2.0550 -0.0750 2.3550 0.0750 ;
        RECT 1.9425 -0.0750 2.0550 0.2250 ;
        RECT 1.6350 -0.0750 1.9425 0.0750 ;
        RECT 1.5150 -0.0750 1.6350 0.1800 ;
        RECT 0.7950 -0.0750 1.5150 0.0750 ;
        RECT 0.6750 -0.0750 0.7950 0.2550 ;
        RECT 0.0000 -0.0750 0.6750 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 2.4750 0.9750 2.7300 1.1250 ;
        RECT 2.3550 0.8700 2.4750 1.1250 ;
        RECT 2.0550 0.9750 2.3550 1.1250 ;
        RECT 1.9425 0.8325 2.0550 1.1250 ;
        RECT 1.6200 0.9750 1.9425 1.1250 ;
        RECT 1.5300 0.8400 1.6200 1.1250 ;
        RECT 0.0000 0.9750 1.5300 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 2.5950 0.2400 2.6550 0.3000 ;
        RECT 2.5950 0.7650 2.6550 0.8250 ;
        RECT 2.4900 0.4950 2.5500 0.5550 ;
        RECT 2.3850 0.1200 2.4450 0.1800 ;
        RECT 2.3850 0.8700 2.4450 0.9300 ;
        RECT 2.2800 0.4950 2.3400 0.5550 ;
        RECT 2.1750 0.2325 2.2350 0.2925 ;
        RECT 2.1750 0.7650 2.2350 0.8250 ;
        RECT 2.0700 0.4950 2.1300 0.5550 ;
        RECT 1.9650 0.1425 2.0250 0.2025 ;
        RECT 1.9650 0.8625 2.0250 0.9225 ;
        RECT 1.8600 0.4950 1.9200 0.5550 ;
        RECT 1.7550 0.1725 1.8150 0.2325 ;
        RECT 1.7550 0.8325 1.8150 0.8925 ;
        RECT 1.6500 0.4950 1.7100 0.5550 ;
        RECT 1.5450 0.1200 1.6050 0.1800 ;
        RECT 1.5450 0.8700 1.6050 0.9300 ;
        RECT 1.4400 0.4950 1.5000 0.5550 ;
        RECT 1.3350 0.2400 1.3950 0.3000 ;
        RECT 1.3350 0.8325 1.3950 0.8925 ;
        RECT 1.2225 0.4950 1.2825 0.5550 ;
        RECT 1.1250 0.6750 1.1850 0.7350 ;
        RECT 1.0200 0.4950 1.0800 0.5550 ;
        RECT 0.9150 0.8325 0.9750 0.8925 ;
        RECT 0.8100 0.4950 0.8700 0.5550 ;
        RECT 0.7050 0.1875 0.7650 0.2475 ;
        RECT 0.7050 0.6825 0.7650 0.7425 ;
        RECT 0.6000 0.4950 0.6600 0.5550 ;
        RECT 0.4950 0.8325 0.5550 0.8925 ;
        RECT 0.3900 0.4950 0.4500 0.5550 ;
        RECT 0.2850 0.6825 0.3450 0.7425 ;
        RECT 0.1875 0.4800 0.2475 0.5400 ;
        RECT 0.0750 0.2100 0.1350 0.2700 ;
        RECT 0.0750 0.8175 0.1350 0.8775 ;
        LAYER M1 ;
        RECT 2.5875 0.2100 2.6625 0.3300 ;
        RECT 2.4675 0.4050 2.6625 0.6150 ;
        RECT 2.5875 0.6900 2.6625 0.8625 ;
        RECT 2.3925 0.2550 2.5875 0.3300 ;
        RECT 2.3175 0.6900 2.5875 0.7950 ;
        RECT 2.3175 0.2550 2.3925 0.5850 ;
        RECT 1.7175 0.4950 2.3175 0.5850 ;
        RECT 2.1675 0.1800 2.2425 0.4200 ;
        RECT 2.1675 0.6675 2.2425 0.8550 ;
        RECT 1.8675 0.3000 2.1675 0.4200 ;
        RECT 1.8675 0.6675 2.1675 0.7575 ;
        RECT 1.7925 0.1500 1.8675 0.4200 ;
        RECT 1.7925 0.6675 1.8675 0.9000 ;
        RECT 1.7325 0.1500 1.7925 0.2550 ;
        RECT 1.7250 0.8250 1.7925 0.9000 ;
        RECT 1.6425 0.3300 1.7175 0.7350 ;
        RECT 1.5675 0.2550 1.6425 0.4050 ;
        RECT 1.0275 0.6600 1.6425 0.7350 ;
        RECT 1.4025 0.2550 1.5675 0.3300 ;
        RECT 1.4925 0.4800 1.5675 0.5850 ;
        RECT 1.3575 0.4050 1.4925 0.5850 ;
        RECT 1.1625 0.8175 1.4250 0.9000 ;
        RECT 1.3275 0.2100 1.4025 0.3300 ;
        RECT 1.2300 0.4650 1.2825 0.5850 ;
        RECT 1.1550 0.2175 1.2300 0.5850 ;
        RECT 0.1575 0.8250 1.1625 0.9000 ;
        RECT 0.9750 0.3450 1.0800 0.5850 ;
        RECT 0.9750 0.6600 1.0275 0.7500 ;
        RECT 0.4725 0.3450 0.9750 0.4200 ;
        RECT 0.2925 0.6750 0.9750 0.7500 ;
        RECT 0.5475 0.4950 0.9000 0.6000 ;
        RECT 0.3675 0.3450 0.4725 0.5850 ;
        RECT 0.2175 0.1800 0.2925 0.5700 ;
        RECT 0.2250 0.6450 0.2925 0.7500 ;
        RECT 0.1125 0.6450 0.2250 0.7200 ;
        RECT 0.1875 0.4500 0.2175 0.5700 ;
        RECT 0.0525 0.7950 0.1575 0.9000 ;
        RECT 0.1125 0.1800 0.1350 0.3000 ;
        RECT 0.0375 0.1800 0.1125 0.7200 ;
        LAYER VIA1 ;
        RECT 2.3625 0.7125 2.4375 0.7875 ;
        RECT 1.2375 0.8175 1.3125 0.8925 ;
        LAYER M2 ;
        RECT 2.3625 0.7125 2.4825 0.7875 ;
        RECT 2.2800 0.7125 2.3625 0.9375 ;
        RECT 1.6125 0.8625 2.2800 0.9375 ;
        RECT 1.5225 0.8175 1.6125 0.9375 ;
        RECT 1.1625 0.8175 1.5225 0.8925 ;
    END
END AO31_0111


MACRO AO31_1000
    CLASS CORE ;
    FOREIGN AO31_1000 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.2600 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 1.1475 0.1500 1.2225 0.9000 ;
        RECT 1.1175 0.1500 1.1475 0.3825 ;
        RECT 1.1175 0.6675 1.1475 0.9000 ;
        END
    END Z
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.8475 0.1125 1.1925 0.1875 ;
        RECT 0.7725 0.1125 0.8475 0.5250 ;
        RECT 0.6525 0.1125 0.7725 0.1875 ;
        VIA 0.8100 0.4425 VIA12_square ;
        END
    END B
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.0675 0.2625 0.5325 0.3375 ;
        VIA 0.2550 0.3000 VIA12_square ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.4725 0.8625 0.9225 0.9375 ;
        RECT 0.3675 0.4350 0.4725 0.9375 ;
        VIA 0.4200 0.5175 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.6525 0.7125 1.0875 0.7875 ;
        RECT 0.5775 0.3975 0.6525 0.7875 ;
        VIA 0.6150 0.5175 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.0050 -0.0750 1.2600 0.0750 ;
        RECT 0.8850 -0.0750 1.0050 0.1800 ;
        RECT 0.1425 -0.0750 0.8850 0.0750 ;
        RECT 0.0675 -0.0750 0.1425 0.2550 ;
        RECT 0.0000 -0.0750 0.0675 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.0050 0.9750 1.2600 1.1250 ;
        RECT 0.9000 0.8250 1.0050 1.1250 ;
        RECT 0.0000 0.9750 0.9000 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.1250 0.1800 1.1850 0.2400 ;
        RECT 1.1250 0.8100 1.1850 0.8700 ;
        RECT 1.0125 0.4950 1.0725 0.5550 ;
        RECT 0.9150 0.1200 0.9750 0.1800 ;
        RECT 0.9150 0.8550 0.9750 0.9150 ;
        RECT 0.8100 0.4800 0.8700 0.5400 ;
        RECT 0.7050 0.2100 0.7650 0.2700 ;
        RECT 0.7050 0.8325 0.7650 0.8925 ;
        RECT 0.5925 0.4950 0.6525 0.5550 ;
        RECT 0.4950 0.6825 0.5550 0.7425 ;
        RECT 0.3900 0.4875 0.4500 0.5475 ;
        RECT 0.2850 0.8325 0.3450 0.8925 ;
        RECT 0.1800 0.4950 0.2400 0.5550 ;
        RECT 0.0750 0.1575 0.1350 0.2175 ;
        RECT 0.0750 0.8100 0.1350 0.8700 ;
        LAYER M1 ;
        RECT 1.0425 0.4650 1.0725 0.5850 ;
        RECT 0.9675 0.2550 1.0425 0.7500 ;
        RECT 0.7725 0.2550 0.9675 0.3300 ;
        RECT 0.1500 0.6750 0.9675 0.7500 ;
        RECT 0.7275 0.4050 0.8925 0.6000 ;
        RECT 0.2550 0.8250 0.7950 0.9000 ;
        RECT 0.6975 0.1800 0.7725 0.3300 ;
        RECT 0.6225 0.4275 0.6525 0.6000 ;
        RECT 0.5475 0.2175 0.6225 0.6000 ;
        RECT 0.3675 0.2175 0.4725 0.6000 ;
        RECT 0.2175 0.2175 0.2925 0.5850 ;
        RECT 0.1725 0.4650 0.2175 0.5850 ;
        RECT 0.0450 0.6750 0.1500 0.9000 ;
    END
END AO31_1000


MACRO AO31_1010
    CLASS CORE ;
    FOREIGN AO31_1010 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.2600 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 1.1475 0.2175 1.2225 0.8325 ;
        RECT 1.1175 0.2175 1.1475 0.3825 ;
        RECT 1.1175 0.6675 1.1475 0.8325 ;
        END
    END Z
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.8475 0.1125 1.1925 0.1875 ;
        RECT 0.7725 0.1125 0.8475 0.5250 ;
        RECT 0.6525 0.1125 0.7725 0.1875 ;
        VIA 0.8100 0.4425 VIA12_square ;
        END
    END B
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.0675 0.2625 0.5325 0.3375 ;
        VIA 0.2550 0.3000 VIA12_square ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.4725 0.8625 0.9225 0.9375 ;
        RECT 0.3675 0.4350 0.4725 0.9375 ;
        VIA 0.4200 0.5175 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.6525 0.7125 1.0875 0.7875 ;
        RECT 0.5775 0.3975 0.6525 0.7875 ;
        VIA 0.6150 0.5175 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.0050 -0.0750 1.2600 0.0750 ;
        RECT 0.8850 -0.0750 1.0050 0.1800 ;
        RECT 0.1425 -0.0750 0.8850 0.0750 ;
        RECT 0.0675 -0.0750 0.1425 0.3225 ;
        RECT 0.0000 -0.0750 0.0675 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.0050 0.9750 1.2600 1.1250 ;
        RECT 0.9000 0.8400 1.0050 1.1250 ;
        RECT 0.0000 0.9750 0.9000 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.1250 0.2700 1.1850 0.3300 ;
        RECT 1.1250 0.7275 1.1850 0.7875 ;
        RECT 1.0125 0.4950 1.0725 0.5550 ;
        RECT 0.9150 0.1200 0.9750 0.1800 ;
        RECT 0.9150 0.8700 0.9750 0.9300 ;
        RECT 0.8100 0.4800 0.8700 0.5400 ;
        RECT 0.7050 0.2400 0.7650 0.3000 ;
        RECT 0.7050 0.8325 0.7650 0.8925 ;
        RECT 0.5925 0.4950 0.6525 0.5550 ;
        RECT 0.4950 0.6825 0.5550 0.7425 ;
        RECT 0.3900 0.4875 0.4500 0.5475 ;
        RECT 0.2850 0.8325 0.3450 0.8925 ;
        RECT 0.1800 0.4950 0.2400 0.5550 ;
        RECT 0.0750 0.2250 0.1350 0.2850 ;
        RECT 0.0750 0.7575 0.1350 0.8175 ;
        LAYER M1 ;
        RECT 1.0425 0.4650 1.0725 0.5850 ;
        RECT 0.9675 0.2550 1.0425 0.7500 ;
        RECT 0.7725 0.2550 0.9675 0.3300 ;
        RECT 0.1425 0.6750 0.9675 0.7500 ;
        RECT 0.7275 0.4050 0.8925 0.6000 ;
        RECT 0.2550 0.8250 0.7950 0.9000 ;
        RECT 0.6975 0.2100 0.7725 0.3300 ;
        RECT 0.6225 0.4275 0.6525 0.6000 ;
        RECT 0.5475 0.2175 0.6225 0.6000 ;
        RECT 0.3675 0.2175 0.4725 0.6000 ;
        RECT 0.2175 0.2175 0.2925 0.5850 ;
        RECT 0.1725 0.4650 0.2175 0.5850 ;
        RECT 0.0675 0.6750 0.1425 0.8475 ;
    END
END AO31_1010


MACRO AO32_0011
    CLASS CORE ;
    FOREIGN AO32_0011 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.8900 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.2775 0.2175 0.3525 0.3675 ;
        RECT 0.2775 0.6675 0.3525 0.8550 ;
        RECT 0.1125 0.2925 0.2775 0.3675 ;
        RECT 0.1125 0.6675 0.2775 0.7425 ;
        RECT 0.0375 0.2925 0.1125 0.7425 ;
        END
    END Z
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.3575 0.4125 1.8225 0.4875 ;
        VIA 1.6800 0.4500 VIA12_square ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.3575 0.2625 1.8225 0.3375 ;
        VIA 1.5150 0.3000 VIA12_square ;
        END
    END B1
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.7425 0.4125 0.8175 0.5925 ;
        RECT 0.2775 0.4125 0.7425 0.4875 ;
        VIA 0.7800 0.5100 VIA12_square ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.9675 0.3900 1.0425 0.9375 ;
        RECT 0.9150 0.3900 0.9675 0.4950 ;
        RECT 0.5175 0.8625 0.9675 0.9375 ;
        VIA 1.0050 0.5325 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.2375 0.8625 1.8225 0.9375 ;
        RECT 1.1625 0.3900 1.2375 0.9375 ;
        VIA 1.2000 0.5175 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.8450 -0.0750 1.8900 0.0750 ;
        RECT 1.7250 -0.0750 1.8450 0.2625 ;
        RECT 0.7875 -0.0750 1.7250 0.0750 ;
        RECT 0.6825 -0.0750 0.7875 0.2400 ;
        RECT 0.5775 -0.0750 0.6825 0.0750 ;
        RECT 0.4725 -0.0750 0.5775 0.2400 ;
        RECT 0.1650 -0.0750 0.4725 0.0750 ;
        RECT 0.0450 -0.0750 0.1650 0.2175 ;
        RECT 0.0000 -0.0750 0.0450 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.6350 0.9750 1.8900 1.1250 ;
        RECT 1.5150 0.8550 1.6350 1.1250 ;
        RECT 0.5850 0.9750 1.5150 1.1250 ;
        RECT 0.4650 0.8250 0.5850 1.1250 ;
        RECT 0.1650 0.9750 0.4650 1.1250 ;
        RECT 0.0450 0.8175 0.1650 1.1250 ;
        RECT 0.0000 0.9750 0.0450 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.7550 0.1725 1.8150 0.2325 ;
        RECT 1.7550 0.7425 1.8150 0.8025 ;
        RECT 1.6500 0.4950 1.7100 0.5550 ;
        RECT 1.5450 0.8550 1.6050 0.9150 ;
        RECT 1.4400 0.4875 1.5000 0.5475 ;
        RECT 1.3350 0.1800 1.3950 0.2400 ;
        RECT 1.3350 0.8325 1.3950 0.8925 ;
        RECT 1.2300 0.4875 1.2900 0.5475 ;
        RECT 1.1250 0.6825 1.1850 0.7425 ;
        RECT 1.0200 0.4650 1.0800 0.5250 ;
        RECT 0.9150 0.8325 0.9750 0.8925 ;
        RECT 0.8025 0.5025 0.8625 0.5625 ;
        RECT 0.7050 0.1575 0.7650 0.2175 ;
        RECT 0.7050 0.6825 0.7650 0.7425 ;
        RECT 0.4950 0.1575 0.5550 0.2175 ;
        RECT 0.4950 0.8325 0.5550 0.8925 ;
        RECT 0.3900 0.4950 0.4500 0.5550 ;
        RECT 0.2850 0.2550 0.3450 0.3150 ;
        RECT 0.2850 0.7650 0.3450 0.8250 ;
        RECT 0.1875 0.4950 0.2475 0.5550 ;
        RECT 0.0750 0.1575 0.1350 0.2175 ;
        RECT 0.0750 0.8325 0.1350 0.8925 ;
        LAYER M1 ;
        RECT 1.7400 0.7050 1.8300 0.8325 ;
        RECT 1.6425 0.3675 1.7925 0.5925 ;
        RECT 1.4400 0.7050 1.7400 0.7800 ;
        RECT 1.6200 0.4875 1.6425 0.5925 ;
        RECT 1.5450 0.2175 1.5675 0.4050 ;
        RECT 1.4700 0.2175 1.5450 0.6300 ;
        RECT 1.4400 0.3300 1.4700 0.6300 ;
        RECT 1.3650 0.7050 1.4400 0.9000 ;
        RECT 1.2900 0.1500 1.3950 0.2700 ;
        RECT 1.1625 0.4350 1.3650 0.6000 ;
        RECT 0.8850 0.8250 1.3650 0.9000 ;
        RECT 0.9375 0.1500 1.2900 0.2250 ;
        RECT 0.5025 0.6750 1.2150 0.7500 ;
        RECT 1.0875 0.3000 1.1175 0.3750 ;
        RECT 1.0125 0.3000 1.0875 0.6000 ;
        RECT 0.9375 0.4650 1.0125 0.6000 ;
        RECT 0.8625 0.1500 0.9375 0.3900 ;
        RECT 0.5025 0.3150 0.8625 0.3900 ;
        RECT 0.5775 0.4725 0.8625 0.6000 ;
        RECT 0.4275 0.3150 0.5025 0.7500 ;
        RECT 0.1875 0.4650 0.4275 0.5850 ;
    END
END AO32_0011


MACRO AO32_0111
    CLASS CORE ;
    FOREIGN AO32_0111 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.3600 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 2.6775 0.2400 2.9925 0.7500 ;
        VIA 2.8350 0.3225 VIA12_slot ;
        VIA 2.8350 0.6675 VIA12_slot ;
        END
    END Z
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.7425 0.2625 0.8175 0.5775 ;
        RECT 0.4275 0.2625 0.7425 0.3375 ;
        RECT 0.3525 0.2625 0.4275 0.4875 ;
        RECT 0.1425 0.4125 0.3525 0.4875 ;
        VIA 0.7800 0.4950 VIA12_square ;
        VIA 0.2250 0.4500 VIA12_square ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.5250 0.4425 0.6300 0.7875 ;
        RECT 0.1500 0.7125 0.5250 0.7875 ;
        VIA 0.5775 0.5250 VIA12_square ;
        END
    END B1
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 2.0325 0.1125 2.1225 0.5775 ;
        RECT 1.1925 0.1125 2.0325 0.1875 ;
        RECT 1.1175 0.1125 1.1925 0.5775 ;
        RECT 1.0575 0.4125 1.1175 0.5775 ;
        VIA 2.0775 0.4950 VIA12_square ;
        VIA 1.1100 0.4950 VIA12_square ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.8075 0.3825 1.9125 0.9375 ;
        RECT 1.2825 0.8625 1.8075 0.9375 ;
        VIA 1.8600 0.4725 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.5375 0.3600 1.6125 0.7875 ;
        RECT 1.0725 0.7125 1.5375 0.7875 ;
        VIA 1.5750 0.5250 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 3.2925 -0.0750 3.3600 0.0750 ;
        RECT 3.2175 -0.0750 3.2925 0.3150 ;
        RECT 2.8950 -0.0750 3.2175 0.0750 ;
        RECT 2.7750 -0.0750 2.8950 0.1950 ;
        RECT 2.4750 -0.0750 2.7750 0.0750 ;
        RECT 2.3550 -0.0750 2.4750 0.2175 ;
        RECT 2.2650 -0.0750 2.3550 0.0750 ;
        RECT 2.1450 -0.0750 2.2650 0.2175 ;
        RECT 1.0050 -0.0750 2.1450 0.0750 ;
        RECT 0.8850 -0.0750 1.0050 0.1875 ;
        RECT 0.1575 -0.0750 0.8850 0.0750 ;
        RECT 0.0525 -0.0750 0.1575 0.2850 ;
        RECT 0.0000 -0.0750 0.0525 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 3.2925 0.9750 3.3600 1.1250 ;
        RECT 3.2175 0.6375 3.2925 1.1250 ;
        RECT 2.8875 0.9750 3.2175 1.1250 ;
        RECT 2.7825 0.7950 2.8875 1.1250 ;
        RECT 2.4750 0.9750 2.7825 1.1250 ;
        RECT 2.3700 0.8025 2.4750 1.1250 ;
        RECT 0.7950 0.9750 2.3700 1.1250 ;
        RECT 0.6750 0.8625 0.7950 1.1250 ;
        RECT 0.3750 0.9750 0.6750 1.1250 ;
        RECT 0.2550 0.8625 0.3750 1.1250 ;
        RECT 0.0000 0.9750 0.2550 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 3.2250 0.2250 3.2850 0.2850 ;
        RECT 3.2250 0.6675 3.2850 0.7275 ;
        RECT 3.2250 0.8325 3.2850 0.8925 ;
        RECT 3.1200 0.4650 3.1800 0.5250 ;
        RECT 3.0150 0.2250 3.0750 0.2850 ;
        RECT 3.0150 0.7575 3.0750 0.8175 ;
        RECT 2.9100 0.4650 2.9700 0.5250 ;
        RECT 2.8050 0.1275 2.8650 0.1875 ;
        RECT 2.8050 0.8250 2.8650 0.8850 ;
        RECT 2.7000 0.4650 2.7600 0.5250 ;
        RECT 2.5950 0.2250 2.6550 0.2850 ;
        RECT 2.5950 0.7575 2.6550 0.8175 ;
        RECT 2.4900 0.4650 2.5500 0.5250 ;
        RECT 2.3850 0.1575 2.4450 0.2175 ;
        RECT 2.3850 0.8325 2.4450 0.8925 ;
        RECT 2.1750 0.1575 2.2350 0.2175 ;
        RECT 2.1750 0.8100 2.2350 0.8700 ;
        RECT 2.0700 0.4725 2.1300 0.5325 ;
        RECT 1.9650 0.6600 2.0250 0.7200 ;
        RECT 1.8600 0.4650 1.9200 0.5250 ;
        RECT 1.7550 0.8100 1.8150 0.8700 ;
        RECT 1.6500 0.4875 1.7100 0.5475 ;
        RECT 1.5450 0.1725 1.6050 0.2325 ;
        RECT 1.5450 0.6600 1.6050 0.7200 ;
        RECT 1.4400 0.4875 1.5000 0.5475 ;
        RECT 1.3350 0.8100 1.3950 0.8700 ;
        RECT 1.2300 0.4650 1.2900 0.5250 ;
        RECT 1.1250 0.6600 1.1850 0.7200 ;
        RECT 1.0200 0.4650 1.0800 0.5250 ;
        RECT 0.9150 0.1200 0.9750 0.1800 ;
        RECT 0.9150 0.7575 0.9750 0.8175 ;
        RECT 0.8100 0.4650 0.8700 0.5250 ;
        RECT 0.7050 0.8700 0.7650 0.9300 ;
        RECT 0.6000 0.4875 0.6600 0.5475 ;
        RECT 0.4950 0.2700 0.5550 0.3300 ;
        RECT 0.4950 0.7200 0.5550 0.7800 ;
        RECT 0.3900 0.4875 0.4500 0.5475 ;
        RECT 0.2850 0.8700 0.3450 0.9300 ;
        RECT 0.1800 0.4650 0.2400 0.5250 ;
        RECT 0.0750 0.2025 0.1350 0.2625 ;
        RECT 0.0750 0.7425 0.1350 0.8025 ;
        LAYER M1 ;
        RECT 2.4900 0.4425 3.2100 0.5475 ;
        RECT 2.9925 0.1950 3.0975 0.3675 ;
        RECT 3.0075 0.6225 3.0825 0.8700 ;
        RECT 2.6625 0.6225 3.0075 0.7125 ;
        RECT 2.6775 0.2775 2.9925 0.3675 ;
        RECT 2.5725 0.1950 2.6775 0.3675 ;
        RECT 2.5875 0.6225 2.6625 0.8700 ;
        RECT 2.4150 0.2925 2.4900 0.7275 ;
        RECT 2.0700 0.2925 2.4150 0.3675 ;
        RECT 1.0875 0.6525 2.4150 0.7275 ;
        RECT 2.0025 0.4425 2.3025 0.5475 ;
        RECT 0.9825 0.8025 2.2650 0.8775 ;
        RECT 1.9950 0.1650 2.0700 0.3675 ;
        RECT 1.1550 0.1650 1.9950 0.2400 ;
        RECT 1.8150 0.3225 1.9200 0.5550 ;
        RECT 1.3350 0.3225 1.8150 0.3975 ;
        RECT 1.4100 0.4725 1.7400 0.5775 ;
        RECT 1.2300 0.3225 1.3350 0.5550 ;
        RECT 1.0800 0.1650 1.1550 0.3375 ;
        RECT 0.9600 0.4125 1.1550 0.5775 ;
        RECT 0.4650 0.2625 1.0800 0.3375 ;
        RECT 0.9075 0.7125 0.9825 0.8775 ;
        RECT 0.1425 0.7125 0.9075 0.7875 ;
        RECT 0.7425 0.4125 0.8850 0.6375 ;
        RECT 0.3825 0.4575 0.6675 0.5775 ;
        RECT 0.1125 0.3900 0.3075 0.5550 ;
        RECT 0.0675 0.7125 0.1425 0.8325 ;
    END
END AO32_0111


MACRO AO32_1000
    CLASS CORE ;
    FOREIGN AO32_1000 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.6800 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1125 0.1500 0.1425 0.3825 ;
        RECT 0.1125 0.6675 0.1425 0.9000 ;
        RECT 0.0375 0.1500 0.1125 0.9000 ;
        END
    END Z
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.1475 0.4125 1.6125 0.4875 ;
        VIA 1.4700 0.4500 VIA12_square ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.1475 0.2625 1.6125 0.3375 ;
        VIA 1.3050 0.3000 VIA12_square ;
        END
    END B1
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.5325 0.4125 0.6075 0.5925 ;
        RECT 0.0675 0.4125 0.5325 0.4875 ;
        VIA 0.5700 0.5100 VIA12_square ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.7575 0.3900 0.8325 0.9375 ;
        RECT 0.7050 0.3900 0.7575 0.4950 ;
        RECT 0.3075 0.8625 0.7575 0.9375 ;
        VIA 0.7950 0.5325 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.0275 0.8625 1.6125 0.9375 ;
        RECT 0.9525 0.3900 1.0275 0.9375 ;
        VIA 0.9900 0.5175 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.6350 -0.0750 1.6800 0.0750 ;
        RECT 1.5150 -0.0750 1.6350 0.2625 ;
        RECT 0.5775 -0.0750 1.5150 0.0750 ;
        RECT 0.4725 -0.0750 0.5775 0.2400 ;
        RECT 0.3675 -0.0750 0.4725 0.0750 ;
        RECT 0.2625 -0.0750 0.3675 0.2400 ;
        RECT 0.0000 -0.0750 0.2625 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.4250 0.9750 1.6800 1.1250 ;
        RECT 1.3050 0.8550 1.4250 1.1250 ;
        RECT 0.3750 0.9750 1.3050 1.1250 ;
        RECT 0.2550 0.8250 0.3750 1.1250 ;
        RECT 0.0000 0.9750 0.2550 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.5450 0.1725 1.6050 0.2325 ;
        RECT 1.5450 0.8100 1.6050 0.8700 ;
        RECT 1.4400 0.4950 1.5000 0.5550 ;
        RECT 1.3350 0.8550 1.3950 0.9150 ;
        RECT 1.2300 0.4875 1.2900 0.5475 ;
        RECT 1.1250 0.1800 1.1850 0.2400 ;
        RECT 1.1250 0.8325 1.1850 0.8925 ;
        RECT 1.0200 0.4875 1.0800 0.5475 ;
        RECT 0.9150 0.6825 0.9750 0.7425 ;
        RECT 0.8100 0.4650 0.8700 0.5250 ;
        RECT 0.7050 0.8325 0.7650 0.8925 ;
        RECT 0.5925 0.5025 0.6525 0.5625 ;
        RECT 0.4950 0.1575 0.5550 0.2175 ;
        RECT 0.4950 0.8100 0.5550 0.8700 ;
        RECT 0.2850 0.1575 0.3450 0.2175 ;
        RECT 0.2850 0.8325 0.3450 0.8925 ;
        RECT 0.1875 0.4875 0.2475 0.5475 ;
        RECT 0.0750 0.1800 0.1350 0.2400 ;
        RECT 0.0750 0.8100 0.1350 0.8700 ;
        LAYER M1 ;
        RECT 1.5225 0.7050 1.6275 0.9000 ;
        RECT 1.4325 0.3675 1.5825 0.5925 ;
        RECT 1.2300 0.7050 1.5225 0.7800 ;
        RECT 1.4100 0.4875 1.4325 0.5925 ;
        RECT 1.3350 0.2175 1.3575 0.4050 ;
        RECT 1.2600 0.2175 1.3350 0.6300 ;
        RECT 1.2300 0.3300 1.2600 0.6300 ;
        RECT 1.1550 0.7050 1.2300 0.9000 ;
        RECT 1.0800 0.1500 1.1850 0.2700 ;
        RECT 0.9525 0.4350 1.1550 0.6000 ;
        RECT 0.6750 0.8250 1.1550 0.9000 ;
        RECT 0.7275 0.1500 1.0800 0.2250 ;
        RECT 0.5700 0.6750 1.0050 0.7500 ;
        RECT 0.8775 0.3000 0.9075 0.3750 ;
        RECT 0.8025 0.3000 0.8775 0.6000 ;
        RECT 0.7275 0.4650 0.8025 0.6000 ;
        RECT 0.6525 0.1500 0.7275 0.3900 ;
        RECT 0.2925 0.3150 0.6525 0.3900 ;
        RECT 0.3675 0.4725 0.6525 0.6000 ;
        RECT 0.4650 0.6750 0.5700 0.9000 ;
        RECT 0.2925 0.6750 0.4650 0.7500 ;
        RECT 0.2175 0.3150 0.2925 0.7500 ;
        RECT 0.1875 0.4575 0.2175 0.5775 ;
    END
END AO32_1000


MACRO AO32_1010
    CLASS CORE ;
    FOREIGN AO32_1010 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.6800 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1125 0.2175 0.1425 0.3825 ;
        RECT 0.1125 0.6675 0.1425 0.8325 ;
        RECT 0.0375 0.2175 0.1125 0.8325 ;
        END
    END Z
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.1475 0.4125 1.6125 0.4875 ;
        VIA 1.4700 0.4500 VIA12_square ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.1475 0.2625 1.6125 0.3375 ;
        VIA 1.3050 0.3000 VIA12_square ;
        END
    END B1
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.5325 0.4125 0.6075 0.5925 ;
        RECT 0.0675 0.4125 0.5325 0.4875 ;
        VIA 0.5700 0.5100 VIA12_square ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.7575 0.3900 0.8325 0.9375 ;
        RECT 0.7050 0.3900 0.7575 0.4950 ;
        RECT 0.3075 0.8625 0.7575 0.9375 ;
        VIA 0.7950 0.5325 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.0275 0.8625 1.6125 0.9375 ;
        RECT 0.9525 0.3900 1.0275 0.9375 ;
        VIA 0.9900 0.5175 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.6350 -0.0750 1.6800 0.0750 ;
        RECT 1.5150 -0.0750 1.6350 0.2625 ;
        RECT 0.5775 -0.0750 1.5150 0.0750 ;
        RECT 0.4725 -0.0750 0.5775 0.2400 ;
        RECT 0.3675 -0.0750 0.4725 0.0750 ;
        RECT 0.2625 -0.0750 0.3675 0.2400 ;
        RECT 0.0000 -0.0750 0.2625 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.4250 0.9750 1.6800 1.1250 ;
        RECT 1.3050 0.8550 1.4250 1.1250 ;
        RECT 0.3750 0.9750 1.3050 1.1250 ;
        RECT 0.2550 0.8250 0.3750 1.1250 ;
        RECT 0.0000 0.9750 0.2550 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.5450 0.1725 1.6050 0.2325 ;
        RECT 1.5450 0.7425 1.6050 0.8025 ;
        RECT 1.4400 0.4950 1.5000 0.5550 ;
        RECT 1.3350 0.8550 1.3950 0.9150 ;
        RECT 1.2300 0.4875 1.2900 0.5475 ;
        RECT 1.1250 0.1800 1.1850 0.2400 ;
        RECT 1.1250 0.8325 1.1850 0.8925 ;
        RECT 1.0200 0.4875 1.0800 0.5475 ;
        RECT 0.9150 0.6825 0.9750 0.7425 ;
        RECT 0.8100 0.4650 0.8700 0.5250 ;
        RECT 0.7050 0.8325 0.7650 0.8925 ;
        RECT 0.5925 0.5025 0.6525 0.5625 ;
        RECT 0.4950 0.1575 0.5550 0.2175 ;
        RECT 0.4950 0.6825 0.5550 0.7425 ;
        RECT 0.2850 0.1575 0.3450 0.2175 ;
        RECT 0.2850 0.8325 0.3450 0.8925 ;
        RECT 0.1875 0.4875 0.2475 0.5475 ;
        RECT 0.0750 0.2700 0.1350 0.3300 ;
        RECT 0.0750 0.7200 0.1350 0.7800 ;
        LAYER M1 ;
        RECT 1.5300 0.7050 1.6200 0.8325 ;
        RECT 1.4325 0.3675 1.5825 0.5925 ;
        RECT 1.2300 0.7050 1.5300 0.7800 ;
        RECT 1.4100 0.4875 1.4325 0.5925 ;
        RECT 1.3350 0.2175 1.3575 0.4050 ;
        RECT 1.2600 0.2175 1.3350 0.6300 ;
        RECT 1.2300 0.3300 1.2600 0.6300 ;
        RECT 1.1550 0.7050 1.2300 0.9000 ;
        RECT 1.0800 0.1500 1.1850 0.2700 ;
        RECT 0.9525 0.4350 1.1550 0.6000 ;
        RECT 0.6750 0.8250 1.1550 0.9000 ;
        RECT 0.7275 0.1500 1.0800 0.2250 ;
        RECT 0.2925 0.6750 1.0050 0.7500 ;
        RECT 0.8775 0.3000 0.9075 0.3750 ;
        RECT 0.8025 0.3000 0.8775 0.6000 ;
        RECT 0.7275 0.4650 0.8025 0.6000 ;
        RECT 0.6525 0.1500 0.7275 0.3900 ;
        RECT 0.2925 0.3150 0.6525 0.3900 ;
        RECT 0.3675 0.4725 0.6525 0.6000 ;
        RECT 0.2175 0.3150 0.2925 0.7500 ;
        RECT 0.1875 0.4575 0.2175 0.5775 ;
    END
END AO32_1010


MACRO AO33_0011
    CLASS CORE ;
    FOREIGN AO33_0011 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.8900 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 1.7775 0.3075 1.8525 0.7425 ;
        RECT 1.6125 0.3075 1.7775 0.3825 ;
        RECT 1.6125 0.6675 1.7775 0.7425 ;
        RECT 1.5375 0.2175 1.6125 0.3825 ;
        RECT 1.5375 0.6675 1.6125 0.8550 ;
        END
    END Z
    PIN B3
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.1550 0.1125 1.6200 0.1875 ;
        RECT 1.1550 0.4125 1.3125 0.4875 ;
        RECT 1.0800 0.1125 1.1550 0.4875 ;
        VIA 1.2300 0.4500 VIA12_square ;
        END
    END B3
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.9300 0.1125 1.0050 0.4200 ;
        RECT 0.4650 0.1125 0.9300 0.1875 ;
        RECT 0.9000 0.3150 0.9300 0.4200 ;
        VIA 0.9675 0.3375 VIA12_square ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.8175 0.5625 1.3200 0.6375 ;
        RECT 0.7125 0.4275 0.8175 0.6375 ;
        VIA 0.7650 0.5025 VIA12_square ;
        END
    END B1
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1500 0.4650 0.2400 0.5850 ;
        RECT 0.1425 0.3675 0.1500 0.5850 ;
        RECT 0.0375 0.3675 0.1425 0.6825 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.4500 0.2625 0.7650 0.3375 ;
        RECT 0.3750 0.2625 0.4500 0.7875 ;
        RECT 0.0600 0.7125 0.3750 0.7875 ;
        VIA 0.4125 0.3600 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.6000 0.4275 0.6300 0.5925 ;
        RECT 0.5250 0.4275 0.6000 0.9375 ;
        RECT 0.0600 0.8625 0.5250 0.9375 ;
        VIA 0.5700 0.5100 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.8450 -0.0750 1.8900 0.0750 ;
        RECT 1.7250 -0.0750 1.8450 0.2175 ;
        RECT 1.4250 -0.0750 1.7250 0.0750 ;
        RECT 1.3050 -0.0750 1.4250 0.1800 ;
        RECT 0.1650 -0.0750 1.3050 0.0750 ;
        RECT 0.0450 -0.0750 0.1650 0.2625 ;
        RECT 0.0000 -0.0750 0.0450 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.8450 0.9750 1.8900 1.1250 ;
        RECT 1.7250 0.8175 1.8450 1.1250 ;
        RECT 1.4250 0.9750 1.7250 1.1250 ;
        RECT 1.3050 0.8700 1.4250 1.1250 ;
        RECT 1.0200 0.9750 1.3050 1.1250 ;
        RECT 0.9150 0.8250 1.0200 1.1250 ;
        RECT 0.0000 0.9750 0.9150 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.7550 0.1575 1.8150 0.2175 ;
        RECT 1.7550 0.8325 1.8150 0.8925 ;
        RECT 1.6425 0.4950 1.7025 0.5550 ;
        RECT 1.5450 0.2775 1.6050 0.3375 ;
        RECT 1.5450 0.7650 1.6050 0.8250 ;
        RECT 1.4400 0.4950 1.5000 0.5550 ;
        RECT 1.3350 0.1200 1.3950 0.1800 ;
        RECT 1.3350 0.8700 1.3950 0.9300 ;
        RECT 1.2300 0.4725 1.2900 0.5325 ;
        RECT 1.1250 0.7500 1.1850 0.8100 ;
        RECT 1.0125 0.4725 1.0725 0.5325 ;
        RECT 0.9150 0.8550 0.9750 0.9150 ;
        RECT 0.8025 0.4950 0.8625 0.5550 ;
        RECT 0.7050 0.1575 0.7650 0.2175 ;
        RECT 0.7050 0.6750 0.7650 0.7350 ;
        RECT 0.5925 0.4725 0.6525 0.5325 ;
        RECT 0.4950 0.8250 0.5550 0.8850 ;
        RECT 0.3900 0.4800 0.4500 0.5400 ;
        RECT 0.2850 0.6750 0.3450 0.7350 ;
        RECT 0.1800 0.4950 0.2400 0.5550 ;
        RECT 0.0750 0.1725 0.1350 0.2325 ;
        RECT 0.0750 0.8025 0.1350 0.8625 ;
        LAYER M1 ;
        RECT 1.4625 0.4650 1.7025 0.5850 ;
        RECT 1.3875 0.2550 1.4625 0.7950 ;
        RECT 1.2300 0.2550 1.3875 0.3300 ;
        RECT 1.2975 0.7125 1.3875 0.7950 ;
        RECT 1.1475 0.4050 1.3125 0.6000 ;
        RECT 1.1550 0.1500 1.2300 0.3300 ;
        RECT 1.1025 0.6750 1.1925 0.8400 ;
        RECT 0.6750 0.1500 1.1550 0.2250 ;
        RECT 1.0050 0.6750 1.1025 0.7500 ;
        RECT 0.9975 0.3000 1.0725 0.5625 ;
        RECT 0.9300 0.6675 1.0050 0.7500 ;
        RECT 0.8775 0.3000 0.9975 0.4050 ;
        RECT 0.2550 0.6675 0.9300 0.7425 ;
        RECT 0.8025 0.4800 0.9225 0.5850 ;
        RECT 0.1500 0.8175 0.8100 0.8925 ;
        RECT 0.7275 0.3300 0.8025 0.5850 ;
        RECT 0.5325 0.3150 0.6525 0.5925 ;
        RECT 0.3225 0.2325 0.4575 0.5850 ;
        RECT 0.0450 0.7725 0.1500 0.8925 ;
        LAYER VIA1 ;
        RECT 1.3425 0.7200 1.4175 0.7950 ;
        RECT 0.6900 0.8175 0.7650 0.8925 ;
        LAYER M2 ;
        RECT 1.3200 0.7200 1.4625 0.7950 ;
        RECT 1.2450 0.7200 1.3200 0.9375 ;
        RECT 0.7800 0.8625 1.2450 0.9375 ;
        RECT 0.6750 0.7725 0.7800 0.9375 ;
    END
END AO33_0011


MACRO AO33_0111
    CLASS CORE ;
    FOREIGN AO33_0111 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.7800 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 3.0975 0.2400 3.4125 0.7500 ;
        VIA 3.2550 0.3225 VIA12_slot ;
        VIA 3.2550 0.6675 VIA12_slot ;
        END
    END Z
    PIN B3
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.1625 0.3825 1.2375 0.7950 ;
        RECT 0.4275 0.7050 1.1625 0.7950 ;
        RECT 0.3525 0.4125 0.4275 0.7950 ;
        RECT 0.1425 0.4125 0.3525 0.4875 ;
        VIA 1.2000 0.4950 VIA12_square ;
        VIA 0.2250 0.4500 VIA12_square ;
        END
    END B3
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.2925 0.2625 0.7650 0.3375 ;
        VIA 0.4500 0.3000 VIA12_square ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.8175 0.4125 1.0125 0.4875 ;
        RECT 0.6525 0.4125 0.8175 0.5775 ;
        RECT 0.5475 0.4125 0.6525 0.4875 ;
        VIA 0.7350 0.5250 VIA12_square ;
        END
    END B1
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 2.4525 0.1125 2.5425 0.5775 ;
        RECT 1.6125 0.1125 2.4525 0.1875 ;
        RECT 1.5375 0.1125 1.6125 0.5775 ;
        RECT 1.4775 0.4125 1.5375 0.5775 ;
        VIA 2.4975 0.4950 VIA12_square ;
        VIA 1.5300 0.4950 VIA12_square ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 2.2275 0.3675 2.3325 0.9375 ;
        RECT 1.6950 0.8625 2.2275 0.9375 ;
        VIA 2.2800 0.4500 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.9575 0.4425 2.0325 0.7875 ;
        RECT 1.4850 0.7125 1.9575 0.7875 ;
        VIA 1.9950 0.5250 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 3.7125 -0.0750 3.7800 0.0750 ;
        RECT 3.6375 -0.0750 3.7125 0.3150 ;
        RECT 3.3150 -0.0750 3.6375 0.0750 ;
        RECT 3.1950 -0.0750 3.3150 0.1950 ;
        RECT 2.8950 -0.0750 3.1950 0.0750 ;
        RECT 2.7750 -0.0750 2.8950 0.2175 ;
        RECT 2.6850 -0.0750 2.7750 0.0750 ;
        RECT 2.5650 -0.0750 2.6850 0.2175 ;
        RECT 1.4250 -0.0750 2.5650 0.0750 ;
        RECT 1.3050 -0.0750 1.4250 0.1875 ;
        RECT 0.1650 -0.0750 1.3050 0.0750 ;
        RECT 0.0450 -0.0750 0.1650 0.2775 ;
        RECT 0.0000 -0.0750 0.0450 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 3.7125 0.9750 3.7800 1.1250 ;
        RECT 3.6375 0.6375 3.7125 1.1250 ;
        RECT 3.3075 0.9750 3.6375 1.1250 ;
        RECT 3.2025 0.8025 3.3075 1.1250 ;
        RECT 2.8950 0.9750 3.2025 1.1250 ;
        RECT 2.7900 0.8025 2.8950 1.1250 ;
        RECT 1.2150 0.9750 2.7900 1.1250 ;
        RECT 1.0950 0.8550 1.2150 1.1250 ;
        RECT 0.7950 0.9750 1.0950 1.1250 ;
        RECT 0.6750 0.8475 0.7950 1.1250 ;
        RECT 0.3750 0.9750 0.6750 1.1250 ;
        RECT 0.2550 0.8475 0.3750 1.1250 ;
        RECT 0.0000 0.9750 0.2550 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 3.6450 0.2250 3.7050 0.2850 ;
        RECT 3.6450 0.6675 3.7050 0.7275 ;
        RECT 3.6450 0.8325 3.7050 0.8925 ;
        RECT 3.5400 0.4650 3.6000 0.5250 ;
        RECT 3.4350 0.2250 3.4950 0.2850 ;
        RECT 3.4350 0.7575 3.4950 0.8175 ;
        RECT 3.3300 0.4650 3.3900 0.5250 ;
        RECT 3.2250 0.1275 3.2850 0.1875 ;
        RECT 3.2250 0.8325 3.2850 0.8925 ;
        RECT 3.1200 0.4650 3.1800 0.5250 ;
        RECT 3.0150 0.2250 3.0750 0.2850 ;
        RECT 3.0150 0.7575 3.0750 0.8175 ;
        RECT 2.9100 0.4650 2.9700 0.5250 ;
        RECT 2.8050 0.1575 2.8650 0.2175 ;
        RECT 2.8050 0.8325 2.8650 0.8925 ;
        RECT 2.5950 0.1575 2.6550 0.2175 ;
        RECT 2.5950 0.8100 2.6550 0.8700 ;
        RECT 2.4900 0.4725 2.5500 0.5325 ;
        RECT 2.3850 0.6600 2.4450 0.7200 ;
        RECT 2.2800 0.4650 2.3400 0.5250 ;
        RECT 2.1750 0.8100 2.2350 0.8700 ;
        RECT 2.0700 0.4875 2.1300 0.5475 ;
        RECT 1.9650 0.1725 2.0250 0.2325 ;
        RECT 1.9650 0.6600 2.0250 0.7200 ;
        RECT 1.8600 0.4875 1.9200 0.5475 ;
        RECT 1.7550 0.8100 1.8150 0.8700 ;
        RECT 1.6500 0.4650 1.7100 0.5250 ;
        RECT 1.5450 0.6600 1.6050 0.7200 ;
        RECT 1.4400 0.4650 1.5000 0.5250 ;
        RECT 1.3350 0.1200 1.3950 0.1800 ;
        RECT 1.3350 0.7575 1.3950 0.8175 ;
        RECT 1.2300 0.4650 1.2900 0.5250 ;
        RECT 1.1250 0.8625 1.1850 0.9225 ;
        RECT 1.0200 0.4650 1.0800 0.5250 ;
        RECT 0.9150 0.7050 0.9750 0.7650 ;
        RECT 0.8100 0.4875 0.8700 0.5475 ;
        RECT 0.7050 0.1725 0.7650 0.2325 ;
        RECT 0.7050 0.8550 0.7650 0.9150 ;
        RECT 0.6000 0.4875 0.6600 0.5475 ;
        RECT 0.4950 0.7050 0.5550 0.7650 ;
        RECT 0.3900 0.4650 0.4500 0.5250 ;
        RECT 0.2850 0.8550 0.3450 0.9150 ;
        RECT 0.1800 0.4725 0.2400 0.5325 ;
        RECT 0.0750 0.1950 0.1350 0.2550 ;
        RECT 0.0750 0.7275 0.1350 0.7875 ;
        LAYER M1 ;
        RECT 2.9100 0.4425 3.6300 0.5475 ;
        RECT 3.4125 0.1950 3.5175 0.3675 ;
        RECT 3.4275 0.6225 3.5025 0.8700 ;
        RECT 3.0825 0.6225 3.4275 0.7125 ;
        RECT 3.0975 0.2775 3.4125 0.3675 ;
        RECT 2.9925 0.1950 3.0975 0.3675 ;
        RECT 3.0075 0.6225 3.0825 0.8700 ;
        RECT 2.8350 0.2925 2.9100 0.7275 ;
        RECT 2.4900 0.2925 2.8350 0.3675 ;
        RECT 1.5075 0.6525 2.8350 0.7275 ;
        RECT 2.4225 0.4425 2.7225 0.5475 ;
        RECT 1.4025 0.8025 2.6850 0.8775 ;
        RECT 2.4150 0.1650 2.4900 0.3675 ;
        RECT 1.5750 0.1650 2.4150 0.2400 ;
        RECT 2.2350 0.3225 2.3400 0.5550 ;
        RECT 1.7550 0.3225 2.2350 0.3975 ;
        RECT 1.8300 0.4725 2.1600 0.5775 ;
        RECT 1.6500 0.3225 1.7550 0.5550 ;
        RECT 1.5000 0.1650 1.5750 0.3375 ;
        RECT 1.3800 0.4125 1.5750 0.5775 ;
        RECT 1.2300 0.2625 1.5000 0.3375 ;
        RECT 1.3275 0.6975 1.4025 0.8775 ;
        RECT 0.1425 0.6975 1.3275 0.7725 ;
        RECT 1.1550 0.4125 1.3050 0.6225 ;
        RECT 1.1550 0.1650 1.2300 0.3375 ;
        RECT 0.6675 0.1650 1.1550 0.2400 ;
        RECT 0.9750 0.3225 1.0800 0.5550 ;
        RECT 0.5175 0.3225 0.9750 0.3975 ;
        RECT 0.5700 0.4725 0.9000 0.5775 ;
        RECT 0.4950 0.2175 0.5175 0.3975 ;
        RECT 0.3825 0.2175 0.4950 0.5550 ;
        RECT 0.1050 0.3825 0.3075 0.5475 ;
        RECT 0.0675 0.6975 0.1425 0.8175 ;
    END
END AO33_0111


MACRO AO33_1000
    CLASS CORE ;
    FOREIGN AO33_1000 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.6800 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 1.5675 0.1500 1.6425 0.9000 ;
        RECT 1.5375 0.1500 1.5675 0.3825 ;
        RECT 1.5375 0.6675 1.5675 0.9000 ;
        END
    END Z
    PIN B3
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.1550 0.1125 1.6200 0.1875 ;
        RECT 1.1550 0.4125 1.3125 0.4875 ;
        RECT 1.0800 0.1125 1.1550 0.4875 ;
        VIA 1.2300 0.4500 VIA12_square ;
        END
    END B3
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.9300 0.1125 1.0050 0.4200 ;
        RECT 0.4650 0.1125 0.9300 0.1875 ;
        RECT 0.9000 0.3150 0.9300 0.4200 ;
        VIA 0.9675 0.3375 VIA12_square ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.8175 0.5625 1.3200 0.6375 ;
        RECT 0.7125 0.4275 0.8175 0.6375 ;
        VIA 0.7650 0.5025 VIA12_square ;
        END
    END B1
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1500 0.4650 0.2400 0.5850 ;
        RECT 0.1425 0.3675 0.1500 0.5850 ;
        RECT 0.0375 0.3675 0.1425 0.6825 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.4500 0.2625 0.7650 0.3375 ;
        RECT 0.3750 0.2625 0.4500 0.7875 ;
        RECT 0.0600 0.7125 0.3750 0.7875 ;
        VIA 0.4125 0.3600 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.6000 0.4275 0.6300 0.5925 ;
        RECT 0.5250 0.4275 0.6000 0.9375 ;
        RECT 0.0600 0.8625 0.5250 0.9375 ;
        VIA 0.5700 0.5100 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.4250 -0.0750 1.6800 0.0750 ;
        RECT 1.3050 -0.0750 1.4250 0.1800 ;
        RECT 0.1650 -0.0750 1.3050 0.0750 ;
        RECT 0.0450 -0.0750 0.1650 0.2625 ;
        RECT 0.0000 -0.0750 0.0450 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.4250 0.9750 1.6800 1.1250 ;
        RECT 1.3050 0.8700 1.4250 1.1250 ;
        RECT 1.0200 0.9750 1.3050 1.1250 ;
        RECT 0.9150 0.8250 1.0200 1.1250 ;
        RECT 0.0000 0.9750 0.9150 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.5450 0.1800 1.6050 0.2400 ;
        RECT 1.5450 0.8100 1.6050 0.8700 ;
        RECT 1.4325 0.4875 1.4925 0.5475 ;
        RECT 1.3350 0.1200 1.3950 0.1800 ;
        RECT 1.3350 0.8700 1.3950 0.9300 ;
        RECT 1.2300 0.4725 1.2900 0.5325 ;
        RECT 1.1250 0.7800 1.1850 0.8400 ;
        RECT 1.0125 0.4725 1.0725 0.5325 ;
        RECT 0.9150 0.8550 0.9750 0.9150 ;
        RECT 0.8025 0.4950 0.8625 0.5550 ;
        RECT 0.7050 0.1575 0.7650 0.2175 ;
        RECT 0.7050 0.6750 0.7650 0.7350 ;
        RECT 0.5925 0.4725 0.6525 0.5325 ;
        RECT 0.4950 0.8250 0.5550 0.8850 ;
        RECT 0.3900 0.4800 0.4500 0.5400 ;
        RECT 0.2850 0.6750 0.3450 0.7350 ;
        RECT 0.1800 0.4950 0.2400 0.5550 ;
        RECT 0.0750 0.1725 0.1350 0.2325 ;
        RECT 0.0750 0.8025 0.1350 0.8625 ;
        LAYER M1 ;
        RECT 1.4625 0.4575 1.4925 0.5775 ;
        RECT 1.3875 0.2550 1.4625 0.7950 ;
        RECT 1.2300 0.2550 1.3875 0.3300 ;
        RECT 1.2975 0.7125 1.3875 0.7950 ;
        RECT 1.1475 0.4050 1.3125 0.6000 ;
        RECT 1.1550 0.1500 1.2300 0.3300 ;
        RECT 1.1025 0.6750 1.1925 0.8700 ;
        RECT 0.6750 0.1500 1.1550 0.2250 ;
        RECT 1.0050 0.6750 1.1025 0.7500 ;
        RECT 0.9975 0.3000 1.0725 0.5625 ;
        RECT 0.9300 0.6675 1.0050 0.7500 ;
        RECT 0.8775 0.3000 0.9975 0.4050 ;
        RECT 0.2550 0.6675 0.9300 0.7425 ;
        RECT 0.8025 0.4800 0.9225 0.5850 ;
        RECT 0.1500 0.8175 0.8100 0.8925 ;
        RECT 0.7275 0.3300 0.8025 0.5850 ;
        RECT 0.5325 0.3150 0.6525 0.5925 ;
        RECT 0.3225 0.2325 0.4575 0.5850 ;
        RECT 0.0450 0.7725 0.1500 0.8925 ;
        LAYER VIA1 ;
        RECT 1.3425 0.7200 1.4175 0.7950 ;
        RECT 0.6900 0.8175 0.7650 0.8925 ;
        LAYER M2 ;
        RECT 1.3200 0.7200 1.4625 0.7950 ;
        RECT 1.2450 0.7200 1.3200 0.9375 ;
        RECT 0.7800 0.8625 1.2450 0.9375 ;
        RECT 0.6750 0.7725 0.7800 0.9375 ;
    END
END AO33_1000


MACRO AO33_1010
    CLASS CORE ;
    FOREIGN AO33_1010 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.6800 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 1.5675 0.2175 1.6425 0.8325 ;
        RECT 1.5375 0.2175 1.5675 0.3825 ;
        RECT 1.5375 0.6675 1.5675 0.8325 ;
        END
    END Z
    PIN B3
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.1550 0.1125 1.6200 0.1875 ;
        RECT 1.1550 0.4125 1.3125 0.4875 ;
        RECT 1.0800 0.1125 1.1550 0.4875 ;
        VIA 1.2300 0.4500 VIA12_square ;
        END
    END B3
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.9300 0.1125 1.0050 0.4200 ;
        RECT 0.4650 0.1125 0.9300 0.1875 ;
        RECT 0.9000 0.3150 0.9300 0.4200 ;
        VIA 0.9675 0.3375 VIA12_square ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.8175 0.5625 1.3200 0.6375 ;
        RECT 0.7125 0.4275 0.8175 0.6375 ;
        VIA 0.7650 0.5025 VIA12_square ;
        END
    END B1
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1500 0.4650 0.2400 0.5850 ;
        RECT 0.1425 0.3675 0.1500 0.5850 ;
        RECT 0.0375 0.3675 0.1425 0.6825 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.4500 0.2625 0.7650 0.3375 ;
        RECT 0.3750 0.2625 0.4500 0.7875 ;
        RECT 0.0600 0.7125 0.3750 0.7875 ;
        VIA 0.4125 0.3600 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.6000 0.4275 0.6300 0.5925 ;
        RECT 0.5250 0.4275 0.6000 0.9375 ;
        RECT 0.0600 0.8625 0.5250 0.9375 ;
        VIA 0.5700 0.5100 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.4250 -0.0750 1.6800 0.0750 ;
        RECT 1.3050 -0.0750 1.4250 0.1800 ;
        RECT 0.1650 -0.0750 1.3050 0.0750 ;
        RECT 0.0450 -0.0750 0.1650 0.2625 ;
        RECT 0.0000 -0.0750 0.0450 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.4250 0.9750 1.6800 1.1250 ;
        RECT 1.3050 0.8700 1.4250 1.1250 ;
        RECT 1.0200 0.9750 1.3050 1.1250 ;
        RECT 0.9150 0.8250 1.0200 1.1250 ;
        RECT 0.0000 0.9750 0.9150 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.5450 0.2700 1.6050 0.3300 ;
        RECT 1.5450 0.7200 1.6050 0.7800 ;
        RECT 1.4325 0.4875 1.4925 0.5475 ;
        RECT 1.3350 0.1200 1.3950 0.1800 ;
        RECT 1.3350 0.8700 1.3950 0.9300 ;
        RECT 1.2300 0.4725 1.2900 0.5325 ;
        RECT 1.1250 0.7500 1.1850 0.8100 ;
        RECT 1.0125 0.4725 1.0725 0.5325 ;
        RECT 0.9150 0.8550 0.9750 0.9150 ;
        RECT 0.8025 0.4950 0.8625 0.5550 ;
        RECT 0.7050 0.1575 0.7650 0.2175 ;
        RECT 0.7050 0.6750 0.7650 0.7350 ;
        RECT 0.5925 0.4725 0.6525 0.5325 ;
        RECT 0.4950 0.8250 0.5550 0.8850 ;
        RECT 0.3900 0.4800 0.4500 0.5400 ;
        RECT 0.2850 0.6750 0.3450 0.7350 ;
        RECT 0.1800 0.4950 0.2400 0.5550 ;
        RECT 0.0750 0.1725 0.1350 0.2325 ;
        RECT 0.0750 0.8025 0.1350 0.8625 ;
        LAYER M1 ;
        RECT 1.4625 0.4575 1.4925 0.5775 ;
        RECT 1.3875 0.2550 1.4625 0.7950 ;
        RECT 1.2300 0.2550 1.3875 0.3300 ;
        RECT 1.2975 0.7125 1.3875 0.7950 ;
        RECT 1.1475 0.4050 1.3125 0.6000 ;
        RECT 1.1550 0.1500 1.2300 0.3300 ;
        RECT 1.1025 0.6750 1.1925 0.8400 ;
        RECT 0.6750 0.1500 1.1550 0.2250 ;
        RECT 1.0050 0.6750 1.1025 0.7500 ;
        RECT 0.9975 0.3000 1.0725 0.5625 ;
        RECT 0.9300 0.6675 1.0050 0.7500 ;
        RECT 0.8775 0.3000 0.9975 0.4050 ;
        RECT 0.2550 0.6675 0.9300 0.7425 ;
        RECT 0.8025 0.4800 0.9225 0.5850 ;
        RECT 0.1500 0.8175 0.8100 0.8925 ;
        RECT 0.7275 0.3300 0.8025 0.5850 ;
        RECT 0.5325 0.3150 0.6525 0.5925 ;
        RECT 0.3225 0.2325 0.4575 0.5850 ;
        RECT 0.0450 0.7725 0.1500 0.8925 ;
        LAYER VIA1 ;
        RECT 1.3425 0.7200 1.4175 0.7950 ;
        RECT 0.6900 0.8175 0.7650 0.8925 ;
        LAYER M2 ;
        RECT 1.3200 0.7200 1.4625 0.7950 ;
        RECT 1.2450 0.7200 1.3200 0.9375 ;
        RECT 0.7800 0.8625 1.2450 0.9375 ;
        RECT 0.6750 0.7725 0.7800 0.9375 ;
    END
END AO33_1010


MACRO AOI211_0011
    CLASS CORE ;
    FOREIGN AOI211_0011 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.8900 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 1.0800 0.1125 1.2300 0.2550 ;
        RECT 0.7575 0.1125 1.0800 0.1875 ;
        RECT 0.6825 0.1125 0.7575 0.9375 ;
        RECT 0.2175 0.8625 0.6825 0.9375 ;
        VIA 1.1550 0.2025 VIA12_square ;
        VIA 0.7200 0.2025 VIA12_square ;
        VIA 0.7200 0.7125 VIA12_square ;
        END
    END ZN
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.9825 0.4125 1.4475 0.4875 ;
        VIA 1.3350 0.4500 VIA12_square ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.9075 0.5625 1.7775 0.6375 ;
        VIA 1.6650 0.6000 VIA12_square ;
        VIA 1.0275 0.6000 VIA12_square ;
        END
    END B
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.8175 0.4575 0.8775 0.5775 ;
        RECT 0.7425 0.3150 0.8175 0.5775 ;
        RECT 0.2475 0.3150 0.7425 0.3900 ;
        RECT 0.1425 0.3150 0.2475 0.5550 ;
        RECT 0.0675 0.3150 0.1425 0.6825 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.5325 0.1125 0.6075 0.6000 ;
        RECT 0.0675 0.1125 0.5325 0.1875 ;
        RECT 0.5025 0.4500 0.5325 0.6000 ;
        VIA 0.5550 0.5250 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.8375 -0.0750 1.8900 0.0750 ;
        RECT 1.7325 -0.0750 1.8375 0.3150 ;
        RECT 1.4250 -0.0750 1.7325 0.0750 ;
        RECT 1.3050 -0.0750 1.4250 0.1875 ;
        RECT 0.9825 -0.0750 1.3050 0.0750 ;
        RECT 0.9075 -0.0750 0.9825 0.2775 ;
        RECT 0.1575 -0.0750 0.9075 0.0750 ;
        RECT 0.0525 -0.0750 0.1575 0.2400 ;
        RECT 0.0000 -0.0750 0.0525 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.4250 0.9750 1.8900 1.1250 ;
        RECT 1.3050 0.8625 1.4250 1.1250 ;
        RECT 0.0000 0.9750 1.3050 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.7550 0.2325 1.8150 0.2925 ;
        RECT 1.7550 0.7350 1.8150 0.7950 ;
        RECT 1.6500 0.4800 1.7100 0.5400 ;
        RECT 1.5450 0.2325 1.6050 0.2925 ;
        RECT 1.4400 0.4875 1.5000 0.5475 ;
        RECT 1.3350 0.1275 1.3950 0.1875 ;
        RECT 1.3350 0.8700 1.3950 0.9300 ;
        RECT 1.2300 0.4875 1.2900 0.5475 ;
        RECT 1.1250 0.2325 1.1850 0.2925 ;
        RECT 1.0200 0.4875 1.0800 0.5475 ;
        RECT 0.9150 0.1875 0.9750 0.2475 ;
        RECT 0.9150 0.8325 0.9750 0.8925 ;
        RECT 0.8100 0.4875 0.8700 0.5475 ;
        RECT 0.7050 0.6825 0.7650 0.7425 ;
        RECT 0.6000 0.4950 0.6600 0.5550 ;
        RECT 0.4950 0.1650 0.5550 0.2250 ;
        RECT 0.4950 0.8325 0.5550 0.8925 ;
        RECT 0.3900 0.4950 0.4500 0.5550 ;
        RECT 0.2850 0.6825 0.3450 0.7425 ;
        RECT 0.1800 0.4650 0.2400 0.5250 ;
        RECT 0.0750 0.1575 0.1350 0.2175 ;
        RECT 0.0750 0.8100 0.1350 0.8700 ;
        LAYER M1 ;
        RECT 1.7325 0.7125 1.8375 0.8175 ;
        RECT 1.5825 0.4200 1.7775 0.6375 ;
        RECT 1.2300 0.7125 1.7325 0.7875 ;
        RECT 1.5375 0.2025 1.6125 0.3375 ;
        RECT 1.2300 0.2625 1.5375 0.3375 ;
        RECT 1.2225 0.4125 1.5075 0.5775 ;
        RECT 1.0725 0.1500 1.2300 0.3375 ;
        RECT 1.1550 0.7125 1.2300 0.9000 ;
        RECT 0.1575 0.8250 1.1550 0.9000 ;
        RECT 0.9525 0.4125 1.0800 0.7500 ;
        RECT 0.2550 0.6675 0.8175 0.7500 ;
        RECT 0.4500 0.1500 0.8025 0.2400 ;
        RECT 0.3825 0.4650 0.6675 0.5850 ;
        RECT 0.0525 0.7875 0.1575 0.9000 ;
    END
END AOI211_0011


MACRO AOI211_0100
    CLASS CORE ;
    FOREIGN AOI211_0100 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.2400 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 4.0350 0.2925 4.1925 0.4125 ;
        RECT 4.0350 0.6450 4.1925 0.7650 ;
        RECT 3.7200 0.2925 4.0350 0.7650 ;
        RECT 3.5625 0.2925 3.7200 0.4125 ;
        RECT 3.5625 0.6450 3.7200 0.7650 ;
        VIA 4.0350 0.3525 VIA12_slot ;
        VIA 4.0350 0.7050 VIA12_slot ;
        VIA 3.7200 0.3525 VIA12_slot ;
        VIA 3.7200 0.7050 VIA12_slot ;
        END
    END ZN
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 9.0975 0.3600 9.1725 0.6450 ;
        RECT 9.0075 0.4800 9.0975 0.6450 ;
        RECT 6.6600 0.4800 9.0075 0.5850 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 4.7250 0.5625 5.0850 0.6375 ;
        RECT 4.6200 0.4125 4.7250 0.6375 ;
        VIA 4.6725 0.5250 VIA12_square ;
        END
    END B
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.3225 0.4350 2.5425 0.5625 ;
        RECT 0.1425 0.4050 0.3225 0.5625 ;
        RECT 0.0675 0.4050 0.1425 0.6825 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 2.7450 0.4125 2.8500 0.6000 ;
        RECT 2.3250 0.4125 2.7450 0.4875 ;
        VIA 2.7975 0.5175 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 9.1875 -0.0750 9.2400 0.0750 ;
        RECT 9.0825 -0.0750 9.1875 0.2400 ;
        RECT 8.7750 -0.0750 9.0825 0.0750 ;
        RECT 8.6550 -0.0750 8.7750 0.2175 ;
        RECT 8.3550 -0.0750 8.6550 0.0750 ;
        RECT 8.2350 -0.0750 8.3550 0.2175 ;
        RECT 7.9350 -0.0750 8.2350 0.0750 ;
        RECT 7.8150 -0.0750 7.9350 0.2175 ;
        RECT 7.5150 -0.0750 7.8150 0.0750 ;
        RECT 7.3950 -0.0750 7.5150 0.2175 ;
        RECT 7.0950 -0.0750 7.3950 0.0750 ;
        RECT 6.9750 -0.0750 7.0950 0.2175 ;
        RECT 6.6750 -0.0750 6.9750 0.0750 ;
        RECT 6.5550 -0.0750 6.6750 0.2175 ;
        RECT 6.2550 -0.0750 6.5550 0.0750 ;
        RECT 6.1350 -0.0750 6.2550 0.2175 ;
        RECT 5.8350 -0.0750 6.1350 0.0750 ;
        RECT 5.7150 -0.0750 5.8350 0.2175 ;
        RECT 5.4150 -0.0750 5.7150 0.0750 ;
        RECT 5.2950 -0.0750 5.4150 0.2175 ;
        RECT 4.9950 -0.0750 5.2950 0.0750 ;
        RECT 4.8750 -0.0750 4.9950 0.1800 ;
        RECT 4.5750 -0.0750 4.8750 0.0750 ;
        RECT 4.4550 -0.0750 4.5750 0.2175 ;
        RECT 2.4750 -0.0750 4.4550 0.0750 ;
        RECT 2.3550 -0.0750 2.4750 0.1800 ;
        RECT 2.0550 -0.0750 2.3550 0.0750 ;
        RECT 1.9350 -0.0750 2.0550 0.1800 ;
        RECT 1.6350 -0.0750 1.9350 0.0750 ;
        RECT 1.5150 -0.0750 1.6350 0.1800 ;
        RECT 1.2150 -0.0750 1.5150 0.0750 ;
        RECT 1.0950 -0.0750 1.2150 0.1800 ;
        RECT 0.7950 -0.0750 1.0950 0.0750 ;
        RECT 0.6750 -0.0750 0.7950 0.1800 ;
        RECT 0.3750 -0.0750 0.6750 0.0750 ;
        RECT 0.2550 -0.0750 0.3750 0.1800 ;
        RECT 0.0000 -0.0750 0.2550 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 8.9850 0.9750 9.2400 1.1250 ;
        RECT 8.8650 0.8700 8.9850 1.1250 ;
        RECT 8.5650 0.9750 8.8650 1.1250 ;
        RECT 8.4450 0.8700 8.5650 1.1250 ;
        RECT 8.1450 0.9750 8.4450 1.1250 ;
        RECT 8.0250 0.8700 8.1450 1.1250 ;
        RECT 7.7250 0.9750 8.0250 1.1250 ;
        RECT 7.6050 0.8700 7.7250 1.1250 ;
        RECT 7.3050 0.9750 7.6050 1.1250 ;
        RECT 7.1850 0.8700 7.3050 1.1250 ;
        RECT 6.8850 0.9750 7.1850 1.1250 ;
        RECT 6.7650 0.8700 6.8850 1.1250 ;
        RECT 0.0000 0.9750 6.7650 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 9.1050 0.1575 9.1650 0.2175 ;
        RECT 9.1050 0.7500 9.1650 0.8100 ;
        RECT 9.0000 0.4950 9.0600 0.5550 ;
        RECT 8.8950 0.2400 8.9550 0.3000 ;
        RECT 8.8950 0.8700 8.9550 0.9300 ;
        RECT 8.7900 0.4950 8.8500 0.5550 ;
        RECT 8.6850 0.1575 8.7450 0.2175 ;
        RECT 8.6850 0.7050 8.7450 0.7650 ;
        RECT 8.5800 0.4950 8.6400 0.5550 ;
        RECT 8.4750 0.2400 8.5350 0.3000 ;
        RECT 8.4750 0.8700 8.5350 0.9300 ;
        RECT 8.3700 0.4950 8.4300 0.5550 ;
        RECT 8.2650 0.1575 8.3250 0.2175 ;
        RECT 8.2650 0.6825 8.3250 0.7425 ;
        RECT 8.1600 0.4950 8.2200 0.5550 ;
        RECT 8.0550 0.2400 8.1150 0.3000 ;
        RECT 8.0550 0.8700 8.1150 0.9300 ;
        RECT 7.9500 0.4950 8.0100 0.5550 ;
        RECT 7.8450 0.1575 7.9050 0.2175 ;
        RECT 7.8450 0.6825 7.9050 0.7425 ;
        RECT 7.7400 0.4950 7.8000 0.5550 ;
        RECT 7.6350 0.2400 7.6950 0.3000 ;
        RECT 7.6350 0.8700 7.6950 0.9300 ;
        RECT 7.5300 0.4950 7.5900 0.5550 ;
        RECT 7.4250 0.1575 7.4850 0.2175 ;
        RECT 7.4250 0.6825 7.4850 0.7425 ;
        RECT 7.3200 0.4950 7.3800 0.5550 ;
        RECT 7.2150 0.2400 7.2750 0.3000 ;
        RECT 7.2150 0.8700 7.2750 0.9300 ;
        RECT 7.1100 0.4950 7.1700 0.5550 ;
        RECT 7.0050 0.1575 7.0650 0.2175 ;
        RECT 7.0050 0.6825 7.0650 0.7425 ;
        RECT 6.9000 0.4950 6.9600 0.5550 ;
        RECT 6.7950 0.2400 6.8550 0.3000 ;
        RECT 6.7950 0.8700 6.8550 0.9300 ;
        RECT 6.6900 0.4950 6.7500 0.5550 ;
        RECT 6.5850 0.1575 6.6450 0.2175 ;
        RECT 6.5850 0.6825 6.6450 0.7425 ;
        RECT 6.3750 0.8325 6.4350 0.8925 ;
        RECT 6.2700 0.4950 6.3300 0.5550 ;
        RECT 6.1650 0.1575 6.2250 0.2175 ;
        RECT 6.1650 0.6825 6.2250 0.7425 ;
        RECT 6.0600 0.4950 6.1200 0.5550 ;
        RECT 5.9550 0.2400 6.0150 0.3000 ;
        RECT 5.9550 0.8325 6.0150 0.8925 ;
        RECT 5.8500 0.4950 5.9100 0.5550 ;
        RECT 5.7450 0.1575 5.8050 0.2175 ;
        RECT 5.7450 0.6825 5.8050 0.7425 ;
        RECT 5.6400 0.4950 5.7000 0.5550 ;
        RECT 5.5350 0.2400 5.5950 0.3000 ;
        RECT 5.5350 0.8325 5.5950 0.8925 ;
        RECT 5.4300 0.4950 5.4900 0.5550 ;
        RECT 5.3250 0.1575 5.3850 0.2175 ;
        RECT 5.3250 0.6825 5.3850 0.7425 ;
        RECT 5.2200 0.4950 5.2800 0.5550 ;
        RECT 5.1150 0.2400 5.1750 0.3000 ;
        RECT 5.1150 0.8325 5.1750 0.8925 ;
        RECT 5.0100 0.4950 5.0700 0.5550 ;
        RECT 4.9050 0.1200 4.9650 0.1800 ;
        RECT 4.9050 0.6825 4.9650 0.7425 ;
        RECT 4.8000 0.4950 4.8600 0.5550 ;
        RECT 4.6950 0.2625 4.7550 0.3225 ;
        RECT 4.6950 0.8325 4.7550 0.8925 ;
        RECT 4.5900 0.4950 4.6500 0.5550 ;
        RECT 4.4850 0.1575 4.5450 0.2175 ;
        RECT 4.4850 0.6825 4.5450 0.7425 ;
        RECT 4.3800 0.4950 4.4400 0.5550 ;
        RECT 4.2750 0.1725 4.3350 0.2325 ;
        RECT 4.2750 0.8325 4.3350 0.8925 ;
        RECT 4.1625 0.4950 4.2225 0.5550 ;
        RECT 4.0650 0.3000 4.1250 0.3600 ;
        RECT 4.0650 0.6825 4.1250 0.7425 ;
        RECT 3.9600 0.4950 4.0200 0.5550 ;
        RECT 3.8550 0.1575 3.9150 0.2175 ;
        RECT 3.8550 0.8325 3.9150 0.8925 ;
        RECT 3.7500 0.4950 3.8100 0.5550 ;
        RECT 3.6450 0.3000 3.7050 0.3600 ;
        RECT 3.6450 0.6825 3.7050 0.7425 ;
        RECT 3.5400 0.4950 3.6000 0.5550 ;
        RECT 3.4350 0.1575 3.4950 0.2175 ;
        RECT 3.4350 0.8325 3.4950 0.8925 ;
        RECT 3.3300 0.4950 3.3900 0.5550 ;
        RECT 3.2250 0.3000 3.2850 0.3600 ;
        RECT 3.2250 0.6825 3.2850 0.7425 ;
        RECT 3.1200 0.4950 3.1800 0.5550 ;
        RECT 3.0150 0.1575 3.0750 0.2175 ;
        RECT 3.0150 0.8325 3.0750 0.8925 ;
        RECT 2.9100 0.4950 2.9700 0.5550 ;
        RECT 2.8050 0.3000 2.8650 0.3600 ;
        RECT 2.8050 0.6825 2.8650 0.7425 ;
        RECT 2.7000 0.4950 2.7600 0.5550 ;
        RECT 2.5950 0.2325 2.6550 0.2925 ;
        RECT 2.5950 0.8325 2.6550 0.8925 ;
        RECT 2.4825 0.4650 2.5425 0.5250 ;
        RECT 2.3850 0.1200 2.4450 0.1800 ;
        RECT 2.3850 0.6675 2.4450 0.7275 ;
        RECT 2.2800 0.4650 2.3400 0.5250 ;
        RECT 2.1750 0.2625 2.2350 0.3225 ;
        RECT 2.1750 0.8325 2.2350 0.8925 ;
        RECT 2.0700 0.4650 2.1300 0.5250 ;
        RECT 1.9650 0.1200 2.0250 0.1800 ;
        RECT 1.8600 0.4650 1.9200 0.5250 ;
        RECT 1.7550 0.2625 1.8150 0.3225 ;
        RECT 1.7550 0.8325 1.8150 0.8925 ;
        RECT 1.6500 0.4650 1.7100 0.5250 ;
        RECT 1.5450 0.1200 1.6050 0.1800 ;
        RECT 1.5450 0.6675 1.6050 0.7275 ;
        RECT 1.4400 0.4650 1.5000 0.5250 ;
        RECT 1.3350 0.2625 1.3950 0.3225 ;
        RECT 1.3350 0.8325 1.3950 0.8925 ;
        RECT 1.2300 0.4650 1.2900 0.5250 ;
        RECT 1.1250 0.1200 1.1850 0.1800 ;
        RECT 1.0200 0.4650 1.0800 0.5250 ;
        RECT 0.9150 0.2625 0.9750 0.3225 ;
        RECT 0.9150 0.8325 0.9750 0.8925 ;
        RECT 0.8100 0.4650 0.8700 0.5250 ;
        RECT 0.7050 0.1200 0.7650 0.1800 ;
        RECT 0.7050 0.6675 0.7650 0.7275 ;
        RECT 0.6000 0.4650 0.6600 0.5250 ;
        RECT 0.4950 0.2625 0.5550 0.3225 ;
        RECT 0.4950 0.8325 0.5550 0.8925 ;
        RECT 0.3900 0.4650 0.4500 0.5250 ;
        RECT 0.2850 0.1200 0.3450 0.1800 ;
        RECT 0.2850 0.6675 0.3450 0.7275 ;
        RECT 0.1800 0.4650 0.2400 0.5250 ;
        RECT 0.0750 0.2325 0.1350 0.2925 ;
        RECT 0.0750 0.8175 0.1350 0.8775 ;
        LAYER M1 ;
        RECT 9.0975 0.7200 9.1725 0.8400 ;
        RECT 8.7525 0.7200 9.0975 0.7950 ;
        RECT 8.8875 0.2025 8.9625 0.4050 ;
        RECT 8.5425 0.2925 8.8875 0.4050 ;
        RECT 8.6775 0.6750 8.7525 0.7950 ;
        RECT 4.4400 0.6750 8.6775 0.7500 ;
        RECT 8.4675 0.2025 8.5425 0.4050 ;
        RECT 8.1225 0.2925 8.4675 0.4050 ;
        RECT 8.0475 0.2025 8.1225 0.4050 ;
        RECT 7.7025 0.2925 8.0475 0.4050 ;
        RECT 7.6275 0.2025 7.7025 0.4050 ;
        RECT 7.2825 0.2925 7.6275 0.4050 ;
        RECT 7.2075 0.2025 7.2825 0.4050 ;
        RECT 6.8625 0.2925 7.2075 0.4050 ;
        RECT 6.7875 0.2025 6.8625 0.4050 ;
        RECT 6.0225 0.2925 6.7875 0.4050 ;
        RECT 0.1575 0.8250 6.4800 0.9000 ;
        RECT 4.3500 0.4800 6.3600 0.5850 ;
        RECT 5.9475 0.2025 6.0225 0.4050 ;
        RECT 5.6025 0.2925 5.9475 0.4050 ;
        RECT 5.5275 0.2025 5.6025 0.4050 ;
        RECT 5.1825 0.2925 5.5275 0.4050 ;
        RECT 5.1075 0.2025 5.1825 0.4050 ;
        RECT 4.7625 0.2925 5.1075 0.4050 ;
        RECT 4.6875 0.2025 4.7625 0.4050 ;
        RECT 4.4175 0.3000 4.6875 0.4050 ;
        RECT 4.1775 0.3300 4.4175 0.4050 ;
        RECT 4.2525 0.1500 4.3575 0.2550 ;
        RECT 2.6625 0.1500 4.2525 0.2250 ;
        RECT 2.6550 0.4800 4.2525 0.5850 ;
        RECT 0.2475 0.6600 4.1925 0.7500 ;
        RECT 2.7750 0.3000 4.1775 0.4050 ;
        RECT 2.5875 0.1500 2.6625 0.3300 ;
        RECT 0.1425 0.2550 2.5875 0.3300 ;
        RECT 0.0525 0.7950 0.1575 0.9000 ;
        RECT 0.0675 0.2025 0.1425 0.3300 ;
        LAYER M2 ;
        RECT 4.0650 0.2925 4.1925 0.4125 ;
        RECT 4.0650 0.6450 4.1925 0.7650 ;
        RECT 3.5625 0.2925 3.6900 0.4125 ;
        RECT 3.5625 0.6450 3.6900 0.7650 ;
    END
END AOI211_0100


MACRO AOI211_0111
    CLASS CORE ;
    FOREIGN AOI211_0111 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.7800 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 1.2075 0.2700 1.5225 0.7800 ;
        VIA 1.3650 0.3525 VIA12_slot ;
        VIA 1.3650 0.6975 VIA12_slot ;
        END
    END ZN
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 3.2925 0.4125 3.5700 0.4875 ;
        RECT 3.2175 0.4125 3.2925 0.6375 ;
        RECT 2.9400 0.5625 3.2175 0.6375 ;
        VIA 3.2550 0.5325 VIA12_square ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 2.6625 0.4125 2.9400 0.4875 ;
        RECT 2.5875 0.4125 2.6625 0.6375 ;
        RECT 2.3100 0.5625 2.5875 0.6375 ;
        VIA 2.6250 0.5325 VIA12_square ;
        END
    END B
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.5625 0.4125 0.8400 0.4875 ;
        RECT 0.4875 0.4125 0.5625 0.6375 ;
        RECT 0.2100 0.5625 0.4875 0.6375 ;
        VIA 0.5250 0.5325 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.6575 0.5625 2.1225 0.6375 ;
        VIA 1.7850 0.6000 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 3.5175 -0.0750 3.7800 0.0750 ;
        RECT 3.4125 -0.0750 3.5175 0.2175 ;
        RECT 3.0975 -0.0750 3.4125 0.0750 ;
        RECT 2.9925 -0.0750 3.0975 0.2175 ;
        RECT 2.6775 -0.0750 2.9925 0.0750 ;
        RECT 2.5725 -0.0750 2.6775 0.2175 ;
        RECT 2.2575 -0.0750 2.5725 0.0750 ;
        RECT 2.1525 -0.0750 2.2575 0.2175 ;
        RECT 0.7950 -0.0750 2.1525 0.0750 ;
        RECT 0.6750 -0.0750 0.7950 0.2175 ;
        RECT 0.3750 -0.0750 0.6750 0.0750 ;
        RECT 0.2550 -0.0750 0.3750 0.2175 ;
        RECT 0.0000 -0.0750 0.2550 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 3.5175 0.9750 3.7800 1.1250 ;
        RECT 3.4125 0.8250 3.5175 1.1250 ;
        RECT 3.0975 0.9750 3.4125 1.1250 ;
        RECT 2.9925 0.8250 3.0975 1.1250 ;
        RECT 0.0000 0.9750 2.9925 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 3.6450 0.3075 3.7050 0.3675 ;
        RECT 3.6450 0.6975 3.7050 0.7575 ;
        RECT 3.5400 0.4950 3.6000 0.5550 ;
        RECT 3.4350 0.1350 3.4950 0.1950 ;
        RECT 3.4350 0.8475 3.4950 0.9075 ;
        RECT 3.3300 0.4950 3.3900 0.5550 ;
        RECT 3.2250 0.3225 3.2850 0.3825 ;
        RECT 3.2250 0.6825 3.2850 0.7425 ;
        RECT 3.1200 0.4950 3.1800 0.5550 ;
        RECT 3.0150 0.1350 3.0750 0.1950 ;
        RECT 3.0150 0.8475 3.0750 0.9075 ;
        RECT 2.9100 0.4950 2.9700 0.5550 ;
        RECT 2.8050 0.3225 2.8650 0.3825 ;
        RECT 2.8050 0.6825 2.8650 0.7425 ;
        RECT 2.7000 0.4950 2.7600 0.5550 ;
        RECT 2.5950 0.1350 2.6550 0.1950 ;
        RECT 2.5950 0.8325 2.6550 0.8925 ;
        RECT 2.4900 0.4950 2.5500 0.5550 ;
        RECT 2.3850 0.3225 2.4450 0.3825 ;
        RECT 2.3850 0.6825 2.4450 0.7425 ;
        RECT 2.2800 0.4950 2.3400 0.5550 ;
        RECT 2.1750 0.1350 2.2350 0.1950 ;
        RECT 2.1750 0.8325 2.2350 0.8925 ;
        RECT 2.0700 0.4950 2.1300 0.5550 ;
        RECT 1.9650 0.3075 2.0250 0.3675 ;
        RECT 1.9650 0.6825 2.0250 0.7425 ;
        RECT 1.7550 0.1575 1.8150 0.2175 ;
        RECT 1.7550 0.8325 1.8150 0.8925 ;
        RECT 1.6500 0.4950 1.7100 0.5550 ;
        RECT 1.5450 0.3225 1.6050 0.3825 ;
        RECT 1.5450 0.6675 1.6050 0.7275 ;
        RECT 1.4400 0.4950 1.5000 0.5550 ;
        RECT 1.3350 0.1575 1.3950 0.2175 ;
        RECT 1.3350 0.8325 1.3950 0.8925 ;
        RECT 1.2300 0.4950 1.2900 0.5550 ;
        RECT 1.1250 0.3225 1.1850 0.3825 ;
        RECT 1.1250 0.6675 1.1850 0.7275 ;
        RECT 1.0200 0.4950 1.0800 0.5550 ;
        RECT 0.9150 0.2250 0.9750 0.2850 ;
        RECT 0.9150 0.8325 0.9750 0.8925 ;
        RECT 0.8100 0.4800 0.8700 0.5400 ;
        RECT 0.7050 0.1500 0.7650 0.2100 ;
        RECT 0.7050 0.6675 0.7650 0.7275 ;
        RECT 0.6000 0.4800 0.6600 0.5400 ;
        RECT 0.4950 0.3000 0.5550 0.3600 ;
        RECT 0.4950 0.8325 0.5550 0.8925 ;
        RECT 0.3900 0.4800 0.4500 0.5400 ;
        RECT 0.2850 0.6675 0.3450 0.7275 ;
        RECT 0.1800 0.4800 0.2400 0.5400 ;
        RECT 0.0750 0.2850 0.1350 0.3450 ;
        RECT 0.0750 0.8100 0.1350 0.8700 ;
        RECT 0.2850 0.1500 0.3450 0.2100 ;
        LAYER M1 ;
        RECT 1.1025 0.3000 3.7350 0.4050 ;
        RECT 3.6225 0.6750 3.7275 0.7800 ;
        RECT 2.8725 0.4800 3.6300 0.5850 ;
        RECT 1.9350 0.6750 3.6225 0.7500 ;
        RECT 2.0325 0.4800 2.7900 0.5850 ;
        RECT 0.1575 0.8250 2.6850 0.9000 ;
        RECT 0.9825 0.1500 1.8450 0.2250 ;
        RECT 1.7475 0.4800 1.8225 0.7200 ;
        RECT 0.9900 0.4800 1.7475 0.5700 ;
        RECT 0.2625 0.6450 1.6275 0.7500 ;
        RECT 0.9075 0.1500 0.9825 0.3675 ;
        RECT 0.1575 0.2925 0.9075 0.3675 ;
        RECT 0.1500 0.4500 0.8775 0.5700 ;
        RECT 0.0525 0.2625 0.1575 0.3675 ;
        RECT 0.0525 0.7875 0.1575 0.9000 ;
    END
END AOI211_0111


MACRO AOI211_1000
    CLASS CORE ;
    FOREIGN AOI211_1000 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.0500 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 0.6075 0.2625 0.6975 0.3675 ;
        RECT 0.5325 0.2625 0.6075 0.7875 ;
        RECT 0.4725 0.6225 0.5325 0.7875 ;
        RECT 0.0675 0.7125 0.4725 0.7875 ;
        VIA 0.6150 0.3075 VIA12_square ;
        VIA 0.5100 0.7050 VIA12_square ;
        END
    END ZN
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.9075 0.3675 0.9825 0.6825 ;
        RECT 0.8175 0.4350 0.9075 0.5550 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.8175 0.8625 0.9825 0.9375 ;
        RECT 0.7125 0.7350 0.8175 0.9375 ;
        RECT 0.4125 0.8625 0.7125 0.9375 ;
        VIA 0.7650 0.8175 VIA12_square ;
        END
    END B
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.4275 0.1125 0.6075 0.1875 ;
        RECT 0.3525 0.1125 0.4275 0.5400 ;
        RECT 0.0675 0.1125 0.3525 0.1875 ;
        VIA 0.3900 0.4575 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1425 0.4350 0.2325 0.5625 ;
        RECT 0.0675 0.3675 0.1425 0.6825 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.9975 -0.0750 1.0500 0.0750 ;
        RECT 0.8925 -0.0750 0.9975 0.2400 ;
        RECT 0.5850 -0.0750 0.8925 0.0750 ;
        RECT 0.4650 -0.0750 0.5850 0.1800 ;
        RECT 0.0000 -0.0750 0.4650 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.0125 0.9750 1.0500 1.1250 ;
        RECT 0.9075 0.7875 1.0125 1.1250 ;
        RECT 0.0000 0.9750 0.9075 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 0.9150 0.1575 0.9750 0.2175 ;
        RECT 0.9150 0.8175 0.9750 0.8775 ;
        RECT 0.8175 0.4650 0.8775 0.5250 ;
        RECT 0.7050 0.1800 0.7650 0.2400 ;
        RECT 0.6000 0.4650 0.6600 0.5250 ;
        RECT 0.4950 0.1200 0.5550 0.1800 ;
        RECT 0.4950 0.8325 0.5550 0.8925 ;
        RECT 0.3900 0.4650 0.4500 0.5250 ;
        RECT 0.2850 0.6900 0.3450 0.7500 ;
        RECT 0.1725 0.4650 0.2325 0.5250 ;
        RECT 0.0750 0.1575 0.1350 0.2175 ;
        RECT 0.0750 0.8100 0.1350 0.8700 ;
        LAYER M1 ;
        RECT 0.7425 0.6300 0.8175 0.9000 ;
        RECT 0.6825 0.1500 0.7950 0.3450 ;
        RECT 0.7125 0.4275 0.7425 0.9000 ;
        RECT 0.6675 0.4275 0.7125 0.7050 ;
        RECT 0.3825 0.2700 0.6825 0.3450 ;
        RECT 0.6000 0.4275 0.6675 0.5550 ;
        RECT 0.2475 0.6450 0.5925 0.7500 ;
        RECT 0.1425 0.8250 0.5850 0.9000 ;
        RECT 0.3075 0.4200 0.5250 0.5700 ;
        RECT 0.3075 0.1500 0.3825 0.3450 ;
        RECT 0.1500 0.1500 0.3075 0.2250 ;
        RECT 0.0450 0.1500 0.1500 0.2625 ;
        RECT 0.0675 0.7800 0.1425 0.9000 ;
    END
END AOI211_1000


MACRO AOI211_1010
    CLASS CORE ;
    FOREIGN AOI211_1010 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.2600 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 1.1025 0.2100 1.2075 0.3300 ;
        RECT 0.6675 0.2550 1.1025 0.3300 ;
        RECT 0.5925 0.2550 0.6675 0.7500 ;
        RECT 0.4800 0.2550 0.5925 0.3750 ;
        RECT 0.2550 0.6750 0.5925 0.7500 ;
        END
    END ZN
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.0200 0.4125 1.1850 0.6375 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.7575 0.4125 0.9225 0.6375 ;
        END
    END B
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1425 0.4500 0.2400 0.5700 ;
        RECT 0.0675 0.3675 0.1425 0.6825 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.3900 0.4500 0.4500 0.5700 ;
        RECT 0.3150 0.2175 0.3900 0.5700 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.0050 -0.0750 1.2600 0.0750 ;
        RECT 0.8850 -0.0750 1.0050 0.1800 ;
        RECT 0.1650 -0.0750 0.8850 0.0750 ;
        RECT 0.0450 -0.0750 0.1650 0.2475 ;
        RECT 0.0000 -0.0750 0.0450 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.2150 0.9750 1.2600 1.1250 ;
        RECT 1.0950 0.7575 1.2150 1.1250 ;
        RECT 0.0000 0.9750 1.0950 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.1250 0.2400 1.1850 0.3000 ;
        RECT 1.1250 0.7650 1.1850 0.8250 ;
        RECT 1.0200 0.4800 1.0800 0.5400 ;
        RECT 0.9150 0.1200 0.9750 0.1800 ;
        RECT 0.8100 0.4800 0.8700 0.5400 ;
        RECT 0.7050 0.2625 0.7650 0.3225 ;
        RECT 0.7050 0.8325 0.7650 0.8925 ;
        RECT 0.4950 0.2850 0.5550 0.3450 ;
        RECT 0.4950 0.8325 0.5550 0.8925 ;
        RECT 0.3900 0.4800 0.4500 0.5400 ;
        RECT 0.2850 0.6825 0.3450 0.7425 ;
        RECT 0.1800 0.4800 0.2400 0.5400 ;
        RECT 0.0750 0.1800 0.1350 0.2400 ;
        RECT 0.0750 0.8175 0.1350 0.8775 ;
        LAYER M1 ;
        RECT 0.1575 0.8250 0.7950 0.9000 ;
        RECT 0.0525 0.7950 0.1575 0.9000 ;
    END
END AOI211_1010


MACRO AOI21_0011
    CLASS CORE ;
    FOREIGN AOI21_0011 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.4700 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 1.0425 0.1125 1.1175 0.7950 ;
        RECT 0.3675 0.1125 1.0425 0.1875 ;
        RECT 0.2625 0.1125 0.3675 0.3150 ;
        VIA 1.0800 0.2025 VIA12_square ;
        VIA 1.0800 0.7125 VIA12_square ;
        VIA 0.3150 0.2325 VIA12_square ;
        END
    END ZN
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.2775 0.4125 0.7425 0.4875 ;
        VIA 0.3975 0.4500 VIA12_square ;
        END
    END B
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.8625 0.2625 0.9675 0.3675 ;
        RECT 0.5025 0.2625 0.8625 0.3375 ;
        VIA 0.7275 0.3000 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.8625 0.4575 0.9675 0.6375 ;
        RECT 0.4575 0.5625 0.8625 0.6375 ;
        VIA 0.9150 0.5325 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.4100 -0.0750 1.4700 0.0750 ;
        RECT 1.3350 -0.0750 1.4100 0.3000 ;
        RECT 0.5925 -0.0750 1.3350 0.0750 ;
        RECT 0.4875 -0.0750 0.5925 0.2400 ;
        RECT 0.1425 -0.0750 0.4875 0.0750 ;
        RECT 0.0675 -0.0750 0.1425 0.2925 ;
        RECT 0.0000 -0.0750 0.0675 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.3750 0.9750 1.4700 1.1250 ;
        RECT 0.2550 0.7950 0.3750 1.1250 ;
        RECT 0.0000 0.9750 0.2550 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.3350 0.2100 1.3950 0.2700 ;
        RECT 1.3350 0.7575 1.3950 0.8175 ;
        RECT 1.2300 0.4800 1.2900 0.5400 ;
        RECT 1.1250 0.6825 1.1850 0.7425 ;
        RECT 1.0200 0.4950 1.0800 0.5550 ;
        RECT 0.9150 0.1725 0.9750 0.2325 ;
        RECT 0.9150 0.8325 0.9750 0.8925 ;
        RECT 0.8100 0.4950 0.8700 0.5550 ;
        RECT 0.7050 0.6825 0.7650 0.7425 ;
        RECT 0.6000 0.4800 0.6600 0.5400 ;
        RECT 0.4950 0.1500 0.5550 0.2100 ;
        RECT 0.4950 0.7350 0.5550 0.7950 ;
        RECT 0.3900 0.4725 0.4500 0.5325 ;
        RECT 0.2850 0.2250 0.3450 0.2850 ;
        RECT 0.2850 0.8175 0.3450 0.8775 ;
        RECT 0.1800 0.4725 0.2400 0.5325 ;
        RECT 0.0750 0.1875 0.1350 0.2475 ;
        RECT 0.0750 0.7200 0.1350 0.7800 ;
        LAYER M1 ;
        RECT 1.3350 0.7125 1.4100 0.9000 ;
        RECT 0.5625 0.8250 1.3350 0.9000 ;
        RECT 1.2375 0.4725 1.3200 0.5475 ;
        RECT 1.1625 0.3150 1.2375 0.5475 ;
        RECT 0.8700 0.1500 1.2300 0.2400 ;
        RECT 0.6750 0.6750 1.2300 0.7500 ;
        RECT 0.7650 0.3150 1.1625 0.3900 ;
        RECT 0.8025 0.4650 1.0800 0.6000 ;
        RECT 0.6900 0.2175 0.7650 0.3900 ;
        RECT 0.6750 0.3150 0.6900 0.3900 ;
        RECT 0.6000 0.3150 0.6750 0.5700 ;
        RECT 0.4875 0.6450 0.5625 0.9000 ;
        RECT 0.1500 0.6450 0.4875 0.7200 ;
        RECT 0.1125 0.4125 0.4800 0.5400 ;
        RECT 0.2175 0.1500 0.4125 0.3300 ;
        RECT 0.0675 0.6450 0.1500 0.8175 ;
    END
END AOI21_0011


MACRO AOI21_0100
    CLASS CORE ;
    FOREIGN AOI21_0100 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.1400 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 3.6225 0.3000 3.7800 0.4200 ;
        RECT 3.6225 0.6450 3.7800 0.7650 ;
        RECT 3.3075 0.3000 3.6225 0.7650 ;
        RECT 3.1500 0.3000 3.3075 0.4200 ;
        RECT 3.1500 0.6450 3.3075 0.7650 ;
        VIA 3.6225 0.3600 VIA12_slot ;
        VIA 3.6225 0.7050 VIA12_slot ;
        VIA 3.3075 0.3600 VIA12_slot ;
        VIA 3.3075 0.7050 VIA12_slot ;
        END
    END ZN
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 6.9375 0.4125 7.1025 0.6375 ;
        RECT 4.5600 0.4800 6.9375 0.5850 ;
        END
    END B
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.2025 0.4125 0.6675 0.4875 ;
        VIA 0.3150 0.4500 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 4.4400 0.4125 4.8225 0.4875 ;
        RECT 4.3350 0.4125 4.4400 0.6225 ;
        VIA 4.3875 0.5325 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 7.0725 -0.0750 7.1400 0.0750 ;
        RECT 6.9975 -0.0750 7.0725 0.2625 ;
        RECT 6.6675 -0.0750 6.9975 0.0750 ;
        RECT 6.5625 -0.0750 6.6675 0.2400 ;
        RECT 6.2475 -0.0750 6.5625 0.0750 ;
        RECT 6.1425 -0.0750 6.2475 0.2400 ;
        RECT 5.8275 -0.0750 6.1425 0.0750 ;
        RECT 5.7225 -0.0750 5.8275 0.2400 ;
        RECT 5.4075 -0.0750 5.7225 0.0750 ;
        RECT 5.3025 -0.0750 5.4075 0.2400 ;
        RECT 4.9875 -0.0750 5.3025 0.0750 ;
        RECT 4.8825 -0.0750 4.9875 0.2400 ;
        RECT 4.5750 -0.0750 4.8825 0.0750 ;
        RECT 4.4700 -0.0750 4.5750 0.2475 ;
        RECT 2.4675 -0.0750 4.4700 0.0750 ;
        RECT 2.3625 -0.0750 2.4675 0.2250 ;
        RECT 2.0475 -0.0750 2.3625 0.0750 ;
        RECT 1.9425 -0.0750 2.0475 0.2250 ;
        RECT 1.6275 -0.0750 1.9425 0.0750 ;
        RECT 1.5225 -0.0750 1.6275 0.2250 ;
        RECT 1.2075 -0.0750 1.5225 0.0750 ;
        RECT 1.1025 -0.0750 1.2075 0.2250 ;
        RECT 0.7875 -0.0750 1.1025 0.0750 ;
        RECT 0.6825 -0.0750 0.7875 0.2250 ;
        RECT 0.3750 -0.0750 0.6825 0.0750 ;
        RECT 0.2550 -0.0750 0.3750 0.1875 ;
        RECT 0.0000 -0.0750 0.2550 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 6.8850 0.9750 7.1400 1.1250 ;
        RECT 6.7650 0.8625 6.8850 1.1250 ;
        RECT 6.4650 0.9750 6.7650 1.1250 ;
        RECT 6.3450 0.8175 6.4650 1.1250 ;
        RECT 6.0450 0.9750 6.3450 1.1250 ;
        RECT 5.9250 0.8175 6.0450 1.1250 ;
        RECT 5.6250 0.9750 5.9250 1.1250 ;
        RECT 5.5050 0.8175 5.6250 1.1250 ;
        RECT 5.2050 0.9750 5.5050 1.1250 ;
        RECT 5.0850 0.8175 5.2050 1.1250 ;
        RECT 4.7850 0.9750 5.0850 1.1250 ;
        RECT 4.6650 0.8175 4.7850 1.1250 ;
        RECT 0.0000 0.9750 4.6650 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 7.0050 0.1575 7.0650 0.2175 ;
        RECT 7.0050 0.7650 7.0650 0.8250 ;
        RECT 6.9000 0.4875 6.9600 0.5475 ;
        RECT 6.7950 0.1800 6.8550 0.2400 ;
        RECT 6.7950 0.8625 6.8550 0.9225 ;
        RECT 6.6900 0.4875 6.7500 0.5475 ;
        RECT 6.5850 0.1575 6.6450 0.2175 ;
        RECT 6.5850 0.6750 6.6450 0.7350 ;
        RECT 6.4800 0.4875 6.5400 0.5475 ;
        RECT 6.3750 0.1800 6.4350 0.2400 ;
        RECT 6.3750 0.8475 6.4350 0.9075 ;
        RECT 6.2700 0.4875 6.3300 0.5475 ;
        RECT 6.1650 0.1575 6.2250 0.2175 ;
        RECT 6.1650 0.6750 6.2250 0.7350 ;
        RECT 6.0600 0.4875 6.1200 0.5475 ;
        RECT 5.9550 0.1800 6.0150 0.2400 ;
        RECT 5.9550 0.8475 6.0150 0.9075 ;
        RECT 5.8500 0.4875 5.9100 0.5475 ;
        RECT 5.7450 0.1575 5.8050 0.2175 ;
        RECT 5.7450 0.6750 5.8050 0.7350 ;
        RECT 5.6400 0.4950 5.7000 0.5550 ;
        RECT 5.5350 0.1800 5.5950 0.2400 ;
        RECT 5.5350 0.8475 5.5950 0.9075 ;
        RECT 5.4300 0.4950 5.4900 0.5550 ;
        RECT 5.3250 0.1575 5.3850 0.2175 ;
        RECT 5.3250 0.6750 5.3850 0.7350 ;
        RECT 5.2200 0.4950 5.2800 0.5550 ;
        RECT 5.1150 0.1800 5.1750 0.2400 ;
        RECT 5.1150 0.8475 5.1750 0.9075 ;
        RECT 5.0100 0.4950 5.0700 0.5550 ;
        RECT 4.9050 0.1575 4.9650 0.2175 ;
        RECT 4.9050 0.6750 4.9650 0.7350 ;
        RECT 4.8000 0.4950 4.8600 0.5550 ;
        RECT 4.6950 0.3225 4.7550 0.3825 ;
        RECT 4.6950 0.8475 4.7550 0.9075 ;
        RECT 4.5900 0.4950 4.6500 0.5550 ;
        RECT 4.4850 0.1575 4.5450 0.2175 ;
        RECT 4.4850 0.7725 4.5450 0.8325 ;
        RECT 4.2750 0.1575 4.3350 0.2175 ;
        RECT 4.2750 0.6750 4.3350 0.7350 ;
        RECT 4.1700 0.4950 4.2300 0.5550 ;
        RECT 4.0650 0.3225 4.1250 0.3825 ;
        RECT 4.0650 0.8325 4.1250 0.8925 ;
        RECT 3.9600 0.4950 4.0200 0.5550 ;
        RECT 3.8550 0.1575 3.9150 0.2175 ;
        RECT 3.8550 0.6750 3.9150 0.7350 ;
        RECT 3.7500 0.4950 3.8100 0.5550 ;
        RECT 3.6450 0.3225 3.7050 0.3825 ;
        RECT 3.6450 0.8325 3.7050 0.8925 ;
        RECT 3.5400 0.4950 3.6000 0.5550 ;
        RECT 3.4350 0.1575 3.4950 0.2175 ;
        RECT 3.4350 0.6750 3.4950 0.7350 ;
        RECT 3.3300 0.4950 3.3900 0.5550 ;
        RECT 3.2250 0.3225 3.2850 0.3825 ;
        RECT 3.2250 0.8325 3.2850 0.8925 ;
        RECT 3.1200 0.4950 3.1800 0.5550 ;
        RECT 3.0150 0.1575 3.0750 0.2175 ;
        RECT 3.0150 0.6750 3.0750 0.7350 ;
        RECT 2.9100 0.4950 2.9700 0.5550 ;
        RECT 2.8050 0.3225 2.8650 0.3825 ;
        RECT 2.8050 0.8325 2.8650 0.8925 ;
        RECT 2.7000 0.4950 2.7600 0.5550 ;
        RECT 2.5950 0.2325 2.6550 0.2925 ;
        RECT 2.5950 0.6750 2.6550 0.7350 ;
        RECT 2.4900 0.4950 2.5500 0.5550 ;
        RECT 2.3850 0.1425 2.4450 0.2025 ;
        RECT 2.3850 0.8325 2.4450 0.8925 ;
        RECT 2.2800 0.4950 2.3400 0.5550 ;
        RECT 2.1750 0.3075 2.2350 0.3675 ;
        RECT 2.1750 0.6750 2.2350 0.7350 ;
        RECT 2.0700 0.4950 2.1300 0.5550 ;
        RECT 1.9650 0.1425 2.0250 0.2025 ;
        RECT 1.9650 0.8325 2.0250 0.8925 ;
        RECT 1.8600 0.4950 1.9200 0.5550 ;
        RECT 1.7550 0.3075 1.8150 0.3675 ;
        RECT 1.7550 0.6750 1.8150 0.7350 ;
        RECT 1.6500 0.4950 1.7100 0.5550 ;
        RECT 1.5450 0.1425 1.6050 0.2025 ;
        RECT 1.4400 0.4950 1.5000 0.5550 ;
        RECT 1.3350 0.3075 1.3950 0.3675 ;
        RECT 1.3350 0.6750 1.3950 0.7350 ;
        RECT 1.2300 0.4950 1.2900 0.5550 ;
        RECT 1.1250 0.1425 1.1850 0.2025 ;
        RECT 1.1250 0.8325 1.1850 0.8925 ;
        RECT 1.0200 0.4950 1.0800 0.5550 ;
        RECT 0.9150 0.3075 0.9750 0.3675 ;
        RECT 0.9150 0.6750 0.9750 0.7350 ;
        RECT 0.8100 0.4950 0.8700 0.5550 ;
        RECT 0.7050 0.1425 0.7650 0.2025 ;
        RECT 0.6000 0.4950 0.6600 0.5550 ;
        RECT 0.4950 0.2925 0.5550 0.3525 ;
        RECT 0.4950 0.6750 0.5550 0.7350 ;
        RECT 0.3900 0.4950 0.4500 0.5550 ;
        RECT 0.2850 0.1275 0.3450 0.1875 ;
        RECT 0.2850 0.8325 0.3450 0.8925 ;
        RECT 0.1800 0.4950 0.2400 0.5550 ;
        RECT 0.0750 0.2325 0.1350 0.2925 ;
        RECT 0.0750 0.7350 0.1350 0.7950 ;
        LAYER M1 ;
        RECT 6.9975 0.7125 7.0725 0.8700 ;
        RECT 6.8625 0.7125 6.9975 0.7875 ;
        RECT 6.8475 0.1500 6.8775 0.2700 ;
        RECT 6.7875 0.6675 6.8625 0.7875 ;
        RECT 6.7725 0.1500 6.8475 0.4050 ;
        RECT 4.5525 0.6675 6.7875 0.7425 ;
        RECT 6.4575 0.3225 6.7725 0.4050 ;
        RECT 6.3525 0.1500 6.4575 0.4050 ;
        RECT 6.0375 0.3225 6.3525 0.4050 ;
        RECT 5.9325 0.1500 6.0375 0.4050 ;
        RECT 5.6175 0.3225 5.9325 0.4050 ;
        RECT 5.5125 0.1500 5.6175 0.4050 ;
        RECT 5.1975 0.3225 5.5125 0.4050 ;
        RECT 5.0925 0.1500 5.1975 0.4050 ;
        RECT 2.7750 0.3225 5.0925 0.4050 ;
        RECT 4.4775 0.6675 4.5525 0.9000 ;
        RECT 0.2475 0.8250 4.4775 0.9000 ;
        RECT 2.6700 0.4800 4.4700 0.5850 ;
        RECT 0.1425 0.6600 4.3725 0.7500 ;
        RECT 2.6625 0.1500 4.3650 0.2250 ;
        RECT 2.5875 0.1500 2.6625 0.3750 ;
        RECT 0.5775 0.3000 2.5875 0.3750 ;
        RECT 0.3975 0.4725 2.5725 0.5775 ;
        RECT 0.4725 0.2625 0.5775 0.3750 ;
        RECT 0.1425 0.2625 0.4725 0.3375 ;
        RECT 0.2325 0.4125 0.3975 0.5775 ;
        RECT 0.1350 0.4725 0.2325 0.5775 ;
        RECT 0.0675 0.1875 0.1425 0.3375 ;
        RECT 0.0675 0.6600 0.1425 0.8250 ;
        LAYER M2 ;
        RECT 3.6525 0.3000 3.7800 0.4200 ;
        RECT 3.6525 0.6450 3.7800 0.7650 ;
        RECT 3.1500 0.3000 3.2775 0.4200 ;
        RECT 3.1500 0.6450 3.2775 0.7650 ;
    END
END AOI21_0100


MACRO AOI21_0111
    CLASS CORE ;
    FOREIGN AOI21_0111 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.9400 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 0.9975 0.2700 1.3125 0.7875 ;
        VIA 1.1550 0.3525 VIA12_slot ;
        VIA 1.1550 0.7050 VIA12_slot ;
        END
    END ZN
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 2.4525 0.4125 2.6925 0.4875 ;
        RECT 2.3775 0.4125 2.4525 0.6375 ;
        RECT 2.0475 0.5625 2.3775 0.6375 ;
        VIA 2.4150 0.5325 VIA12_square ;
        END
    END B
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.5625 0.4125 0.8025 0.4875 ;
        RECT 0.4875 0.4125 0.5625 0.6375 ;
        RECT 0.1425 0.5625 0.4875 0.6375 ;
        VIA 0.5250 0.5250 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.8225 0.4125 2.0625 0.4875 ;
        RECT 1.7475 0.4125 1.8225 0.6375 ;
        RECT 1.4325 0.5625 1.7475 0.6375 ;
        VIA 1.7850 0.5325 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 2.8800 -0.0750 2.9400 0.0750 ;
        RECT 2.7900 -0.0750 2.8800 0.3000 ;
        RECT 2.4675 -0.0750 2.7900 0.0750 ;
        RECT 2.3625 -0.0750 2.4675 0.2400 ;
        RECT 2.0550 -0.0750 2.3625 0.0750 ;
        RECT 1.9500 -0.0750 2.0550 0.2475 ;
        RECT 0.7650 -0.0750 1.9500 0.0750 ;
        RECT 0.6600 -0.0750 0.7650 0.2250 ;
        RECT 0.3675 -0.0750 0.6600 0.0750 ;
        RECT 0.2625 -0.0750 0.3675 0.2250 ;
        RECT 0.0000 -0.0750 0.2625 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 2.6850 0.9750 2.9400 1.1250 ;
        RECT 2.5650 0.8175 2.6850 1.1250 ;
        RECT 2.2650 0.9750 2.5650 1.1250 ;
        RECT 2.1450 0.8175 2.2650 1.1250 ;
        RECT 0.0000 0.9750 2.1450 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 2.8050 0.2025 2.8650 0.2625 ;
        RECT 2.8050 0.6975 2.8650 0.7575 ;
        RECT 2.7000 0.4875 2.7600 0.5475 ;
        RECT 2.5950 0.2475 2.6550 0.3075 ;
        RECT 2.5950 0.8475 2.6550 0.9075 ;
        RECT 2.4900 0.4875 2.5500 0.5475 ;
        RECT 2.3850 0.1575 2.4450 0.2175 ;
        RECT 2.3850 0.6750 2.4450 0.7350 ;
        RECT 2.2800 0.4950 2.3400 0.5550 ;
        RECT 2.1750 0.3225 2.2350 0.3825 ;
        RECT 2.1750 0.8475 2.2350 0.9075 ;
        RECT 2.0700 0.4950 2.1300 0.5550 ;
        RECT 1.9650 0.1575 2.0250 0.2175 ;
        RECT 1.9650 0.7725 2.0250 0.8325 ;
        RECT 1.7550 0.1575 1.8150 0.2175 ;
        RECT 1.7550 0.6750 1.8150 0.7350 ;
        RECT 1.6500 0.4950 1.7100 0.5550 ;
        RECT 1.5450 0.3225 1.6050 0.3825 ;
        RECT 1.5450 0.8325 1.6050 0.8925 ;
        RECT 1.4400 0.4950 1.5000 0.5550 ;
        RECT 1.3350 0.1575 1.3950 0.2175 ;
        RECT 1.3350 0.6750 1.3950 0.7350 ;
        RECT 1.2300 0.4950 1.2900 0.5550 ;
        RECT 1.1250 0.3075 1.1850 0.3675 ;
        RECT 1.1250 0.8325 1.1850 0.8925 ;
        RECT 1.0200 0.4950 1.0800 0.5550 ;
        RECT 0.9150 0.1575 0.9750 0.2175 ;
        RECT 0.9150 0.6750 0.9750 0.7350 ;
        RECT 0.8100 0.4950 0.8700 0.5550 ;
        RECT 0.7050 0.1350 0.7650 0.1950 ;
        RECT 0.7050 0.8325 0.7650 0.8925 ;
        RECT 0.6000 0.4950 0.6600 0.5550 ;
        RECT 0.4950 0.3075 0.5550 0.3675 ;
        RECT 0.4950 0.6750 0.5550 0.7350 ;
        RECT 0.3900 0.4950 0.4500 0.5550 ;
        RECT 0.2850 0.1425 0.3450 0.2025 ;
        RECT 0.2850 0.8325 0.3450 0.8925 ;
        RECT 0.1800 0.4950 0.2400 0.5550 ;
        RECT 0.0750 0.2625 0.1350 0.3225 ;
        RECT 0.0750 0.7350 0.1350 0.7950 ;
        LAYER M1 ;
        RECT 2.7825 0.6675 2.8800 0.7950 ;
        RECT 2.0400 0.4800 2.7900 0.5850 ;
        RECT 2.0325 0.6675 2.7825 0.7425 ;
        RECT 2.5875 0.2100 2.6625 0.4050 ;
        RECT 1.2975 0.3225 2.5875 0.4050 ;
        RECT 1.9575 0.6675 2.0325 0.9000 ;
        RECT 0.2475 0.8250 1.9575 0.9000 ;
        RECT 0.9900 0.4800 1.8675 0.5850 ;
        RECT 0.1425 0.6600 1.8525 0.7500 ;
        RECT 0.9150 0.1500 1.8450 0.2250 ;
        RECT 0.9900 0.3000 1.2975 0.4050 ;
        RECT 0.8400 0.1500 0.9150 0.3750 ;
        RECT 0.1575 0.4725 0.8925 0.5775 ;
        RECT 0.1425 0.3000 0.8400 0.3750 ;
        RECT 0.0675 0.2175 0.1425 0.3750 ;
        RECT 0.0675 0.6600 0.1425 0.8250 ;
    END
END AOI21_0111


MACRO AOI21_1000
    CLASS CORE ;
    FOREIGN AOI21_1000 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.0500 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.7350 0.1500 0.7950 0.3825 ;
        RECT 0.6600 0.1500 0.7350 0.7500 ;
        RECT 0.4650 0.1500 0.6600 0.2250 ;
        RECT 0.2550 0.6750 0.6600 0.7500 ;
        END
    END ZN
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.9075 0.3675 0.9825 0.6825 ;
        RECT 0.8100 0.4725 0.9075 0.5925 ;
        END
    END B
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1500 0.4725 0.2700 0.5475 ;
        RECT 0.0450 0.3675 0.1500 0.6825 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.3825 0.3000 0.4575 0.5700 ;
        RECT 0.3525 0.3000 0.3825 0.3825 ;
        RECT 0.2775 0.2175 0.3525 0.3825 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.9900 -0.0750 1.0500 0.0750 ;
        RECT 0.9000 -0.0750 0.9900 0.2475 ;
        RECT 0.1650 -0.0750 0.9000 0.0750 ;
        RECT 0.0450 -0.0750 0.1650 0.2325 ;
        RECT 0.0000 -0.0750 0.0450 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.9825 0.9750 1.0500 1.1250 ;
        RECT 0.9075 0.7875 0.9825 1.1250 ;
        RECT 0.0000 0.9750 0.9075 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 0.9150 0.1575 0.9750 0.2175 ;
        RECT 0.9150 0.8175 0.9750 0.8775 ;
        RECT 0.8100 0.5025 0.8700 0.5625 ;
        RECT 0.7050 0.1575 0.7650 0.2175 ;
        RECT 0.7050 0.8325 0.7650 0.8925 ;
        RECT 0.4950 0.1575 0.5550 0.2175 ;
        RECT 0.4950 0.8325 0.5550 0.8925 ;
        RECT 0.3900 0.4800 0.4500 0.5400 ;
        RECT 0.2850 0.6825 0.3450 0.7425 ;
        RECT 0.1800 0.4800 0.2400 0.5400 ;
        RECT 0.0750 0.1575 0.1350 0.2175 ;
        RECT 0.0750 0.8175 0.1350 0.8775 ;
        LAYER M1 ;
        RECT 0.1575 0.8250 0.7950 0.9000 ;
        RECT 0.0525 0.7950 0.1575 0.9000 ;
    END
END AOI21_1000


MACRO AOI21_1010
    CLASS CORE ;
    FOREIGN AOI21_1010 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.0500 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.7350 0.1500 0.7725 0.3825 ;
        RECT 0.6600 0.1500 0.7350 0.7500 ;
        RECT 0.4650 0.1500 0.6600 0.2250 ;
        RECT 0.2550 0.6750 0.6600 0.7500 ;
        END
    END ZN
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.9075 0.3675 0.9825 0.6825 ;
        RECT 0.8100 0.4500 0.9075 0.5700 ;
        END
    END B
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1500 0.4725 0.2700 0.5475 ;
        RECT 0.0450 0.3675 0.1500 0.6825 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.3825 0.3000 0.4575 0.5700 ;
        RECT 0.3525 0.3000 0.3825 0.3825 ;
        RECT 0.2775 0.2175 0.3525 0.3825 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.9900 -0.0750 1.0500 0.0750 ;
        RECT 0.9000 -0.0750 0.9900 0.2625 ;
        RECT 0.1650 -0.0750 0.9000 0.0750 ;
        RECT 0.0450 -0.0750 0.1650 0.2775 ;
        RECT 0.0000 -0.0750 0.0450 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.9825 0.9750 1.0500 1.1250 ;
        RECT 0.9075 0.7875 0.9825 1.1250 ;
        RECT 0.0000 0.9750 0.9075 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 0.9150 0.1725 0.9750 0.2325 ;
        RECT 0.9150 0.8175 0.9750 0.8775 ;
        RECT 0.8100 0.4800 0.8700 0.5400 ;
        RECT 0.7050 0.2400 0.7650 0.3000 ;
        RECT 0.7050 0.8325 0.7650 0.8925 ;
        RECT 0.4950 0.1575 0.5550 0.2175 ;
        RECT 0.4950 0.8325 0.5550 0.8925 ;
        RECT 0.3900 0.4800 0.4500 0.5400 ;
        RECT 0.2850 0.6825 0.3450 0.7425 ;
        RECT 0.1800 0.4800 0.2400 0.5400 ;
        RECT 0.0750 0.2025 0.1350 0.2625 ;
        RECT 0.0750 0.8175 0.1350 0.8775 ;
        LAYER M1 ;
        RECT 0.1575 0.8250 0.7950 0.9000 ;
        RECT 0.0525 0.7950 0.1575 0.9000 ;
    END
END AOI21_1010


MACRO AOI221_0011
    CLASS CORE ;
    FOREIGN AOI221_0011 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.5200 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 1.3725 0.1650 1.8825 0.2400 ;
        RECT 1.2525 0.1125 1.3725 0.2400 ;
        RECT 0.7275 0.1125 1.2525 0.1875 ;
        RECT 0.7275 0.6225 0.7575 0.7875 ;
        RECT 0.6525 0.1125 0.7275 0.7875 ;
        VIA 1.8000 0.2025 VIA12_square ;
        VIA 1.3650 0.2025 VIA12_square ;
        VIA 0.7050 0.7050 VIA12_square ;
        VIA 0.6900 0.1950 VIA12_square ;
        END
    END ZN
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.4025 0.5625 1.7175 0.6375 ;
        RECT 1.3275 0.4125 1.4025 0.6375 ;
        RECT 1.0125 0.4125 1.3275 0.4875 ;
        VIA 1.3650 0.5100 VIA12_square ;
        END
    END C
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 2.2725 0.3150 2.4525 0.6375 ;
        RECT 1.7625 0.3150 2.2725 0.3900 ;
        RECT 1.6875 0.3150 1.7625 0.5700 ;
        RECT 1.6425 0.4500 1.6875 0.5700 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 2.0325 0.8625 2.3475 0.9375 ;
        RECT 1.9575 0.4125 2.0325 0.9375 ;
        RECT 1.6425 0.4125 1.9575 0.4875 ;
        VIA 1.9950 0.5250 VIA12_square ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.8175 0.4575 0.8775 0.5775 ;
        RECT 0.7425 0.3150 0.8175 0.5775 ;
        RECT 0.2475 0.3150 0.7425 0.3900 ;
        RECT 0.1425 0.3150 0.2475 0.5550 ;
        RECT 0.0675 0.3150 0.1425 0.6825 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.5625 0.8625 1.0275 0.9375 ;
        RECT 0.4875 0.4500 0.5625 0.9375 ;
        RECT 0.4575 0.4500 0.4875 0.6000 ;
        VIA 0.5100 0.5250 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 2.4675 -0.0750 2.5200 0.0750 ;
        RECT 2.3625 -0.0750 2.4675 0.2400 ;
        RECT 1.6125 -0.0750 2.3625 0.0750 ;
        RECT 1.5375 -0.0750 1.6125 0.2775 ;
        RECT 1.1925 -0.0750 1.5375 0.0750 ;
        RECT 1.1175 -0.0750 1.1925 0.2775 ;
        RECT 0.9825 -0.0750 1.1175 0.0750 ;
        RECT 0.9075 -0.0750 0.9825 0.2775 ;
        RECT 0.1575 -0.0750 0.9075 0.0750 ;
        RECT 0.0525 -0.0750 0.1575 0.2400 ;
        RECT 0.0000 -0.0750 0.0525 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 2.2650 0.9750 2.5200 1.1250 ;
        RECT 2.1450 0.8625 2.2650 1.1250 ;
        RECT 1.8450 0.9750 2.1450 1.1250 ;
        RECT 1.7250 0.8250 1.8450 1.1250 ;
        RECT 0.0000 0.9750 1.7250 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 2.3850 0.1575 2.4450 0.2175 ;
        RECT 2.3850 0.7350 2.4450 0.7950 ;
        RECT 2.2800 0.4800 2.3400 0.5400 ;
        RECT 2.1750 0.8700 2.2350 0.9300 ;
        RECT 2.0700 0.4950 2.1300 0.5550 ;
        RECT 1.9650 0.1650 2.0250 0.2250 ;
        RECT 1.9650 0.6975 2.0250 0.7575 ;
        RECT 1.8600 0.4950 1.9200 0.5550 ;
        RECT 1.7550 0.8325 1.8150 0.8925 ;
        RECT 1.6500 0.4800 1.7100 0.5400 ;
        RECT 1.5450 0.1875 1.6050 0.2475 ;
        RECT 1.5450 0.6825 1.6050 0.7425 ;
        RECT 1.4400 0.4800 1.5000 0.5400 ;
        RECT 1.3350 0.2550 1.3950 0.3150 ;
        RECT 1.3350 0.8325 1.3950 0.8925 ;
        RECT 1.2300 0.4800 1.2900 0.5400 ;
        RECT 1.1250 0.1875 1.1850 0.2475 ;
        RECT 1.1250 0.6825 1.1850 0.7425 ;
        RECT 0.9150 0.1875 0.9750 0.2475 ;
        RECT 0.9150 0.8325 0.9750 0.8925 ;
        RECT 0.8100 0.4875 0.8700 0.5475 ;
        RECT 0.7050 0.6825 0.7650 0.7425 ;
        RECT 0.6000 0.4950 0.6600 0.5550 ;
        RECT 0.4950 0.1650 0.5550 0.2250 ;
        RECT 0.4950 0.8325 0.5550 0.8925 ;
        RECT 0.3900 0.4950 0.4500 0.5550 ;
        RECT 0.2850 0.6825 0.3450 0.7425 ;
        RECT 0.1800 0.4650 0.2400 0.5250 ;
        RECT 0.0750 0.1575 0.1350 0.2175 ;
        RECT 0.0750 0.8100 0.1350 0.8700 ;
        LAYER M1 ;
        RECT 2.3625 0.7125 2.4675 0.8175 ;
        RECT 2.0550 0.7125 2.3625 0.7875 ;
        RECT 1.8525 0.4650 2.1375 0.5925 ;
        RECT 1.7175 0.1500 2.0700 0.2400 ;
        RECT 1.9350 0.6750 2.0550 0.7875 ;
        RECT 1.0950 0.6750 1.9350 0.7500 ;
        RECT 1.2000 0.4575 1.5300 0.5625 ;
        RECT 1.2825 0.1500 1.4475 0.3450 ;
        RECT 0.1575 0.8250 1.4250 0.9000 ;
        RECT 0.2550 0.6675 0.9300 0.7500 ;
        RECT 0.4500 0.1500 0.8025 0.2400 ;
        RECT 0.3825 0.4650 0.6675 0.5850 ;
        RECT 0.0525 0.7875 0.1575 0.9000 ;
    END
END AOI221_0011


MACRO AOI221_0111
    CLASS CORE ;
    FOREIGN AOI221_0111 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.5200 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 1.6275 0.2625 1.9425 0.7650 ;
        VIA 1.7850 0.3450 VIA12_slot ;
        VIA 1.7850 0.6825 VIA12_slot ;
        END
    END ZN
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.4100 0.7125 1.4775 0.7875 ;
        RECT 1.2900 0.6000 1.4100 0.7875 ;
        RECT 0.9225 0.7125 1.2900 0.7875 ;
        VIA 1.3500 0.6825 VIA12_square ;
        END
    END C
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.6975 0.4125 0.8025 0.9375 ;
        RECT 0.1575 0.8625 0.6975 0.9375 ;
        VIA 0.7500 0.4875 VIA12_square ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.9525 0.4125 1.4775 0.4875 ;
        VIA 1.0650 0.4500 VIA12_square ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1575 0.4500 0.2325 0.5700 ;
        RECT 0.0525 0.3675 0.1575 0.6825 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.4575 0.1125 0.5625 0.1875 ;
        RECT 0.3525 0.1125 0.4575 0.5700 ;
        RECT 0.0675 0.1125 0.3525 0.1875 ;
        VIA 0.3975 0.4875 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 2.2650 -0.0750 2.5200 0.0750 ;
        RECT 2.1450 -0.0750 2.2650 0.1875 ;
        RECT 1.8450 -0.0750 2.1450 0.0750 ;
        RECT 1.7250 -0.0750 1.8450 0.1950 ;
        RECT 1.4175 -0.0750 1.7250 0.0750 ;
        RECT 1.3125 -0.0750 1.4175 0.2475 ;
        RECT 0.7875 -0.0750 1.3125 0.0750 ;
        RECT 0.6825 -0.0750 0.7875 0.2475 ;
        RECT 0.1650 -0.0750 0.6825 0.0750 ;
        RECT 0.0450 -0.0750 0.1650 0.2175 ;
        RECT 0.0000 -0.0750 0.0450 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 2.2650 0.9750 2.5200 1.1250 ;
        RECT 2.1450 0.8325 2.2650 1.1250 ;
        RECT 1.8375 0.9750 2.1450 1.1250 ;
        RECT 1.7325 0.8250 1.8375 1.1250 ;
        RECT 1.4175 0.9750 1.7325 1.1250 ;
        RECT 1.3125 0.8100 1.4175 1.1250 ;
        RECT 0.0000 0.9750 1.3125 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 2.3850 0.1725 2.4450 0.2325 ;
        RECT 2.3850 0.6900 2.4450 0.7500 ;
        RECT 2.2725 0.4650 2.3325 0.5250 ;
        RECT 2.1750 0.1275 2.2350 0.1875 ;
        RECT 2.1750 0.8400 2.2350 0.9000 ;
        RECT 2.0700 0.4800 2.1300 0.5400 ;
        RECT 1.9650 0.2250 2.0250 0.2850 ;
        RECT 1.9650 0.7200 2.0250 0.7800 ;
        RECT 1.8600 0.4800 1.9200 0.5400 ;
        RECT 1.7550 0.1275 1.8150 0.1875 ;
        RECT 1.7550 0.8475 1.8150 0.9075 ;
        RECT 1.6500 0.4800 1.7100 0.5400 ;
        RECT 1.5450 0.2250 1.6050 0.2850 ;
        RECT 1.5450 0.7200 1.6050 0.7800 ;
        RECT 1.4400 0.4800 1.5000 0.5400 ;
        RECT 1.3350 0.1575 1.3950 0.2175 ;
        RECT 1.3350 0.8325 1.3950 0.8925 ;
        RECT 1.2300 0.4800 1.2900 0.5400 ;
        RECT 1.1250 0.1575 1.1850 0.2175 ;
        RECT 1.1250 0.7350 1.1850 0.7950 ;
        RECT 1.0200 0.4875 1.0800 0.5475 ;
        RECT 0.9150 0.8175 0.9750 0.8775 ;
        RECT 0.8025 0.4650 0.8625 0.5250 ;
        RECT 0.7050 0.1575 0.7650 0.2175 ;
        RECT 0.7050 0.6675 0.7650 0.7275 ;
        RECT 0.4950 0.2175 0.5550 0.2775 ;
        RECT 0.4950 0.8325 0.5550 0.8925 ;
        RECT 0.3900 0.4800 0.4500 0.5400 ;
        RECT 0.2850 0.6900 0.3450 0.7500 ;
        RECT 0.1725 0.4800 0.2325 0.5400 ;
        RECT 0.0750 0.1575 0.1350 0.2175 ;
        RECT 0.0750 0.7950 0.1350 0.8550 ;
        LAYER M1 ;
        RECT 2.4075 0.1500 2.4825 0.7575 ;
        RECT 2.3625 0.1500 2.4075 0.2550 ;
        RECT 2.1825 0.6825 2.4075 0.7575 ;
        RECT 2.2575 0.3300 2.3325 0.5775 ;
        RECT 2.2425 0.3300 2.2575 0.4050 ;
        RECT 2.1075 0.2625 2.2425 0.4050 ;
        RECT 2.1075 0.4800 2.1825 0.7575 ;
        RECT 1.5225 0.4800 2.1075 0.5625 ;
        RECT 1.9425 0.1950 2.0325 0.3825 ;
        RECT 1.9575 0.6375 2.0325 0.8325 ;
        RECT 1.6125 0.6375 1.9575 0.7275 ;
        RECT 1.6275 0.2925 1.9425 0.3825 ;
        RECT 1.5225 0.1950 1.6275 0.3825 ;
        RECT 1.5375 0.6375 1.6125 0.8325 ;
        RECT 1.4175 0.4575 1.5225 0.5625 ;
        RECT 1.3425 0.6375 1.4325 0.7350 ;
        RECT 1.2675 0.3300 1.3425 0.7350 ;
        RECT 1.1925 0.3300 1.2675 0.5700 ;
        RECT 0.8700 0.1500 1.2150 0.2550 ;
        RECT 1.1025 0.6450 1.1925 0.8325 ;
        RECT 0.9375 0.3300 1.1100 0.5700 ;
        RECT 0.7875 0.6450 1.1025 0.7200 ;
        RECT 0.8925 0.7950 0.9975 0.9000 ;
        RECT 0.1575 0.8250 0.8925 0.9000 ;
        RECT 0.6825 0.3300 0.8625 0.5700 ;
        RECT 0.6825 0.6450 0.7875 0.7500 ;
        RECT 0.5325 0.1875 0.6075 0.7200 ;
        RECT 0.4950 0.1875 0.5325 0.3300 ;
        RECT 0.3750 0.6450 0.5325 0.7200 ;
        RECT 0.4200 0.4050 0.4500 0.5700 ;
        RECT 0.3075 0.2175 0.4200 0.5700 ;
        RECT 0.2550 0.6450 0.3750 0.7500 ;
        RECT 0.0525 0.7725 0.1575 0.9000 ;
        LAYER VIA1 ;
        RECT 2.2575 0.4200 2.3325 0.4950 ;
        RECT 1.0125 0.1650 1.0875 0.2400 ;
        RECT 0.5325 0.3075 0.6075 0.3825 ;
        LAYER M2 ;
        RECT 2.1675 0.4200 2.3775 0.4950 ;
        RECT 2.0925 0.1125 2.1675 0.4950 ;
        RECT 1.0875 0.1125 2.0925 0.1875 ;
        RECT 1.0125 0.1125 1.0875 0.3375 ;
        RECT 0.6075 0.2625 1.0125 0.3375 ;
        RECT 0.5325 0.2625 0.6075 0.5625 ;
    END
END AOI221_0111


MACRO AOI221_1000
    CLASS CORE ;
    FOREIGN AOI221_1000 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.4700 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 0.3825 0.4125 0.8475 0.4875 ;
        VIA 0.5625 0.4500 VIA12_square ;
        END
    END ZN
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.8475 0.8625 1.3125 0.9375 ;
        RECT 0.7725 0.5625 0.8475 0.9375 ;
        RECT 0.6225 0.5625 0.7725 0.6375 ;
        VIA 0.7350 0.6000 VIA12_square ;
        END
    END C
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.9675 0.1125 1.0425 0.5850 ;
        RECT 0.4425 0.1125 0.9675 0.1875 ;
        VIA 1.0050 0.5025 VIA12_square ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.3275 0.3675 1.4025 0.6375 ;
        RECT 1.2225 0.4650 1.3275 0.6375 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1575 0.4500 0.2325 0.5700 ;
        RECT 0.0525 0.3675 0.1575 0.6825 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.2475 0.2625 0.7125 0.3375 ;
        VIA 0.3525 0.3000 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.0050 -0.0750 1.4700 0.0750 ;
        RECT 0.8850 -0.0750 1.0050 0.1800 ;
        RECT 0.1650 -0.0750 0.8850 0.0750 ;
        RECT 0.0450 -0.0750 0.1650 0.2175 ;
        RECT 0.0000 -0.0750 0.0450 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.2150 0.9750 1.4700 1.1250 ;
        RECT 1.0950 0.8625 1.2150 1.1250 ;
        RECT 0.0000 0.9750 1.0950 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.3350 0.1575 1.3950 0.2175 ;
        RECT 1.3350 0.8175 1.3950 0.8775 ;
        RECT 1.2300 0.4950 1.2900 0.5550 ;
        RECT 1.1250 0.8625 1.1850 0.9225 ;
        RECT 1.0200 0.4875 1.0800 0.5475 ;
        RECT 0.9150 0.1200 0.9750 0.1800 ;
        RECT 0.9150 0.8175 0.9750 0.8775 ;
        RECT 0.8025 0.4800 0.8625 0.5400 ;
        RECT 0.7050 0.1575 0.7650 0.2175 ;
        RECT 0.7050 0.8175 0.7650 0.8775 ;
        RECT 0.4950 0.1575 0.5550 0.2175 ;
        RECT 0.4950 0.7950 0.5550 0.8550 ;
        RECT 0.3900 0.4800 0.4500 0.5400 ;
        RECT 0.2850 0.6900 0.3450 0.7500 ;
        RECT 0.1725 0.4800 0.2325 0.5400 ;
        RECT 0.0750 0.1575 0.1350 0.2175 ;
        RECT 0.0750 0.7950 0.1350 0.8550 ;
        LAYER M1 ;
        RECT 1.2225 0.1500 1.4250 0.2550 ;
        RECT 1.3125 0.7125 1.4175 0.9000 ;
        RECT 0.9975 0.7125 1.3125 0.7875 ;
        RECT 1.1475 0.1500 1.2225 0.3300 ;
        RECT 0.8100 0.2550 1.1475 0.3300 ;
        RECT 0.9375 0.4050 1.1475 0.6300 ;
        RECT 0.8925 0.7125 0.9975 0.9000 ;
        RECT 0.7875 0.4050 0.8625 0.5700 ;
        RECT 0.7350 0.1500 0.8100 0.3300 ;
        RECT 0.4650 0.7950 0.7950 0.9000 ;
        RECT 0.6825 0.4050 0.7875 0.6825 ;
        RECT 0.6000 0.1500 0.7350 0.2250 ;
        RECT 0.5250 0.1500 0.6000 0.7200 ;
        RECT 0.4650 0.1500 0.5250 0.2550 ;
        RECT 0.3750 0.6450 0.5250 0.7200 ;
        RECT 0.1575 0.8250 0.4650 0.9000 ;
        RECT 0.3900 0.4500 0.4500 0.5700 ;
        RECT 0.3075 0.2175 0.3900 0.5700 ;
        RECT 0.2550 0.6450 0.3750 0.7500 ;
        RECT 0.0525 0.7725 0.1575 0.9000 ;
    END
END AOI221_1000


MACRO AOI221_1010
    CLASS CORE ;
    FOREIGN AOI221_1010 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.4700 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 0.3825 0.4125 0.8475 0.4875 ;
        VIA 0.5625 0.4500 VIA12_square ;
        END
    END ZN
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.8475 0.8625 1.3125 0.9375 ;
        RECT 0.7725 0.5625 0.8475 0.9375 ;
        RECT 0.6225 0.5625 0.7725 0.6375 ;
        VIA 0.7350 0.6000 VIA12_square ;
        END
    END C
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.9675 0.1125 1.0425 0.5850 ;
        RECT 0.4425 0.1125 0.9675 0.1875 ;
        VIA 1.0050 0.5025 VIA12_square ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.3275 0.3675 1.4025 0.6375 ;
        RECT 1.2225 0.4650 1.3275 0.6375 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1575 0.4500 0.2325 0.5700 ;
        RECT 0.0525 0.3675 0.1575 0.6825 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.2475 0.2625 0.7125 0.3375 ;
        VIA 0.3525 0.3000 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.0050 -0.0750 1.4700 0.0750 ;
        RECT 0.8850 -0.0750 1.0050 0.1800 ;
        RECT 0.1650 -0.0750 0.8850 0.0750 ;
        RECT 0.0450 -0.0750 0.1650 0.2175 ;
        RECT 0.0000 -0.0750 0.0450 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.2150 0.9750 1.4700 1.1250 ;
        RECT 1.0950 0.8625 1.2150 1.1250 ;
        RECT 0.0000 0.9750 1.0950 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.3350 0.1575 1.3950 0.2175 ;
        RECT 1.3350 0.8175 1.3950 0.8775 ;
        RECT 1.2300 0.4950 1.2900 0.5550 ;
        RECT 1.1250 0.8625 1.1850 0.9225 ;
        RECT 1.0200 0.4875 1.0800 0.5475 ;
        RECT 0.9150 0.1200 0.9750 0.1800 ;
        RECT 0.9150 0.8175 0.9750 0.8775 ;
        RECT 0.8025 0.4800 0.8625 0.5400 ;
        RECT 0.7050 0.1575 0.7650 0.2175 ;
        RECT 0.7050 0.8175 0.7650 0.8775 ;
        RECT 0.4950 0.1575 0.5550 0.2175 ;
        RECT 0.4950 0.7950 0.5550 0.8550 ;
        RECT 0.3900 0.4800 0.4500 0.5400 ;
        RECT 0.2850 0.6900 0.3450 0.7500 ;
        RECT 0.1725 0.4800 0.2325 0.5400 ;
        RECT 0.0750 0.1575 0.1350 0.2175 ;
        RECT 0.0750 0.7950 0.1350 0.8550 ;
        LAYER M1 ;
        RECT 1.2225 0.1500 1.4250 0.2550 ;
        RECT 1.3125 0.7125 1.4175 0.9000 ;
        RECT 0.9975 0.7125 1.3125 0.7875 ;
        RECT 1.1475 0.1500 1.2225 0.3300 ;
        RECT 0.8100 0.2550 1.1475 0.3300 ;
        RECT 0.9375 0.4050 1.1475 0.6300 ;
        RECT 0.8925 0.7125 0.9975 0.9000 ;
        RECT 0.7875 0.4050 0.8625 0.5700 ;
        RECT 0.7350 0.1500 0.8100 0.3300 ;
        RECT 0.4650 0.7950 0.7950 0.9000 ;
        RECT 0.6825 0.4050 0.7875 0.6825 ;
        RECT 0.6000 0.1500 0.7350 0.2250 ;
        RECT 0.5250 0.1500 0.6000 0.7200 ;
        RECT 0.4650 0.1500 0.5250 0.2550 ;
        RECT 0.3750 0.6450 0.5250 0.7200 ;
        RECT 0.1575 0.8250 0.4650 0.9000 ;
        RECT 0.3900 0.4500 0.4500 0.5700 ;
        RECT 0.3075 0.2175 0.3900 0.5700 ;
        RECT 0.2550 0.6450 0.3750 0.7500 ;
        RECT 0.0525 0.7725 0.1575 0.9000 ;
    END
END AOI221_1010


MACRO AOI222_0011
    CLASS CORE ;
    FOREIGN AOI222_0011 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.9400 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 1.1925 0.2925 1.2825 0.3675 ;
        RECT 1.1175 0.2925 1.1925 0.7875 ;
        RECT 0.7275 0.7125 1.1175 0.7875 ;
        RECT 0.5625 0.6600 0.7275 0.7875 ;
        VIA 1.2000 0.3300 VIA12_square ;
        VIA 0.6450 0.7125 VIA12_square ;
        END
    END ZN
    PIN C2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 2.2875 0.2625 2.7075 0.3375 ;
        RECT 2.2125 0.2625 2.2875 0.4875 ;
        RECT 2.0175 0.4125 2.2125 0.4875 ;
        VIA 2.6250 0.3000 VIA12_square ;
        VIA 2.1150 0.4500 VIA12_square ;
        END
    END C2
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 2.4075 0.4650 2.5125 0.6375 ;
        RECT 2.0175 0.5625 2.4075 0.6375 ;
        VIA 2.4600 0.5400 VIA12_square ;
        END
    END C1
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.7625 0.4425 1.8675 0.6375 ;
        RECT 1.3725 0.5625 1.7625 0.6375 ;
        RECT 1.2675 0.4425 1.3725 0.6375 ;
        VIA 1.8150 0.5175 VIA12_square ;
        VIA 1.3200 0.5250 VIA12_square ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.6275 0.2625 2.0625 0.3375 ;
        RECT 1.5225 0.2625 1.6275 0.4500 ;
        VIA 1.5750 0.3750 VIA12_square ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.9675 0.2625 1.0425 0.5625 ;
        RECT 0.2175 0.2625 0.9675 0.3375 ;
        VIA 1.0050 0.4800 VIA12_square ;
        VIA 0.3000 0.3000 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.3525 0.4125 0.8175 0.4875 ;
        VIA 0.5250 0.4500 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 2.8875 -0.0750 2.9400 0.0750 ;
        RECT 2.7825 -0.0750 2.8875 0.2400 ;
        RECT 2.0550 -0.0750 2.7825 0.0750 ;
        RECT 1.9350 -0.0750 2.0550 0.1800 ;
        RECT 1.2150 -0.0750 1.9350 0.0750 ;
        RECT 1.0950 -0.0750 1.2150 0.2175 ;
        RECT 1.0050 -0.0750 1.0950 0.0750 ;
        RECT 0.8850 -0.0750 1.0050 0.2175 ;
        RECT 0.1425 -0.0750 0.8850 0.0750 ;
        RECT 0.0675 -0.0750 0.1425 0.3075 ;
        RECT 0.0000 -0.0750 0.0675 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 2.6850 0.9750 2.9400 1.1250 ;
        RECT 2.5650 0.8250 2.6850 1.1250 ;
        RECT 2.2650 0.9750 2.5650 1.1250 ;
        RECT 2.1450 0.8250 2.2650 1.1250 ;
        RECT 0.0000 0.9750 2.1450 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 2.8050 0.1575 2.8650 0.2175 ;
        RECT 2.8050 0.6975 2.8650 0.7575 ;
        RECT 2.7000 0.4800 2.7600 0.5400 ;
        RECT 2.5950 0.8325 2.6550 0.8925 ;
        RECT 2.4900 0.4950 2.5500 0.5550 ;
        RECT 2.3850 0.2625 2.4450 0.3225 ;
        RECT 2.3850 0.6825 2.4450 0.7425 ;
        RECT 2.2875 0.4950 2.3475 0.5550 ;
        RECT 2.1750 0.8325 2.2350 0.8925 ;
        RECT 2.0700 0.4800 2.1300 0.5400 ;
        RECT 1.9650 0.1200 2.0250 0.1800 ;
        RECT 1.9650 0.6825 2.0250 0.7425 ;
        RECT 1.8525 0.4800 1.9125 0.5400 ;
        RECT 1.7550 0.8325 1.8150 0.8925 ;
        RECT 1.6425 0.4950 1.7025 0.5550 ;
        RECT 1.5450 0.1575 1.6050 0.2175 ;
        RECT 1.5450 0.6825 1.6050 0.7425 ;
        RECT 1.4475 0.4950 1.5075 0.5550 ;
        RECT 1.3350 0.8325 1.3950 0.8925 ;
        RECT 1.2300 0.4800 1.2900 0.5400 ;
        RECT 1.1250 0.1575 1.1850 0.2175 ;
        RECT 1.1250 0.6825 1.1850 0.7425 ;
        RECT 0.9150 0.1575 0.9750 0.2175 ;
        RECT 0.9150 0.8325 0.9750 0.8925 ;
        RECT 0.8100 0.4650 0.8700 0.5250 ;
        RECT 0.7050 0.6825 0.7650 0.7425 ;
        RECT 0.6000 0.4950 0.6600 0.5550 ;
        RECT 0.4950 0.1575 0.5550 0.2175 ;
        RECT 0.4950 0.8325 0.5550 0.8925 ;
        RECT 0.3900 0.4950 0.4500 0.5550 ;
        RECT 0.2850 0.6825 0.3450 0.7425 ;
        RECT 0.1800 0.4800 0.2400 0.5400 ;
        RECT 0.0750 0.2175 0.1350 0.2775 ;
        RECT 0.0750 0.8100 0.1350 0.8700 ;
        LAYER M1 ;
        RECT 2.7825 0.6750 2.8875 0.7800 ;
        RECT 1.0950 0.6750 2.7825 0.7500 ;
        RECT 2.6925 0.3150 2.7675 0.5700 ;
        RECT 2.6625 0.3150 2.6925 0.3900 ;
        RECT 2.5875 0.2175 2.6625 0.3900 ;
        RECT 2.2875 0.4650 2.5875 0.5925 ;
        RECT 1.8600 0.2550 2.4750 0.3300 ;
        RECT 2.0175 0.4125 2.2125 0.6000 ;
        RECT 1.7775 0.4050 1.9425 0.6000 ;
        RECT 1.7850 0.1500 1.8600 0.3300 ;
        RECT 0.1575 0.8250 1.8450 0.9000 ;
        RECT 1.3950 0.1500 1.7850 0.2250 ;
        RECT 1.6275 0.4650 1.7025 0.5850 ;
        RECT 1.5225 0.3000 1.6275 0.5850 ;
        RECT 1.4475 0.4650 1.5225 0.5850 ;
        RECT 1.2900 0.1500 1.3950 0.3675 ;
        RECT 1.1625 0.4425 1.3725 0.6000 ;
        RECT 0.8100 0.2925 1.2900 0.3675 ;
        RECT 0.7800 0.4425 1.0875 0.5475 ;
        RECT 0.2550 0.6675 0.9000 0.7500 ;
        RECT 0.7350 0.1500 0.8100 0.3675 ;
        RECT 0.4650 0.1500 0.7350 0.2250 ;
        RECT 0.5850 0.4650 0.6600 0.5850 ;
        RECT 0.4725 0.3300 0.5850 0.5850 ;
        RECT 0.3900 0.4650 0.4725 0.5850 ;
        RECT 0.3150 0.2025 0.3600 0.3825 ;
        RECT 0.2400 0.2025 0.3150 0.5550 ;
        RECT 0.1500 0.4725 0.2400 0.5550 ;
        RECT 0.0525 0.7875 0.1575 0.9000 ;
    END
END AOI222_0011


MACRO AOI222_0111
    CLASS CORE ;
    FOREIGN AOI222_0111 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.7300 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 1.8375 0.2625 2.1525 0.7575 ;
        VIA 1.9950 0.3450 VIA12_slot ;
        VIA 1.9950 0.6750 VIA12_slot ;
        END
    END ZN
    PIN C2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.3425 0.4125 1.7025 0.4875 ;
        RECT 1.2375 0.3825 1.3425 0.4875 ;
        VIA 1.4025 0.4500 VIA12_square ;
        END
    END C2
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.1625 0.7125 1.5975 0.7875 ;
        RECT 1.0875 0.4125 1.1625 0.7875 ;
        VIA 1.1250 0.4950 VIA12_square ;
        END
    END C1
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.9525 0.8625 1.4475 0.9375 ;
        RECT 0.8775 0.4350 0.9525 0.9375 ;
        VIA 0.9150 0.5175 VIA12_square ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.6450 0.4125 0.7500 0.9375 ;
        RECT 0.2175 0.8625 0.6450 0.9375 ;
        VIA 0.6975 0.4950 VIA12_square ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1500 0.4425 0.2400 0.5700 ;
        RECT 0.0600 0.3675 0.1500 0.6825 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.4200 0.1125 0.5325 0.1875 ;
        RECT 0.3450 0.1125 0.4200 0.4425 ;
        RECT 0.0675 0.1125 0.3450 0.1875 ;
        VIA 0.3825 0.3600 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 2.4750 -0.0750 2.7300 0.0750 ;
        RECT 2.3550 -0.0750 2.4750 0.1875 ;
        RECT 2.0550 -0.0750 2.3550 0.0750 ;
        RECT 1.9350 -0.0750 2.0550 0.1950 ;
        RECT 1.6125 -0.0750 1.9350 0.0750 ;
        RECT 1.5375 -0.0750 1.6125 0.2475 ;
        RECT 0.9825 -0.0750 1.5375 0.0750 ;
        RECT 0.9075 -0.0750 0.9825 0.2475 ;
        RECT 0.1425 -0.0750 0.9075 0.0750 ;
        RECT 0.0675 -0.0750 0.1425 0.2475 ;
        RECT 0.0000 -0.0750 0.0675 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 2.4750 0.9750 2.7300 1.1250 ;
        RECT 2.3550 0.8325 2.4750 1.1250 ;
        RECT 2.0325 0.9750 2.3550 1.1250 ;
        RECT 1.9575 0.8175 2.0325 1.1250 ;
        RECT 1.6275 0.9750 1.9575 1.1250 ;
        RECT 1.5225 0.6750 1.6275 1.1250 ;
        RECT 1.2150 0.9750 1.5225 1.1250 ;
        RECT 1.1100 0.8025 1.2150 1.1250 ;
        RECT 0.0000 0.9750 1.1100 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 2.5950 0.1725 2.6550 0.2325 ;
        RECT 2.5950 0.6900 2.6550 0.7500 ;
        RECT 2.4825 0.4650 2.5425 0.5250 ;
        RECT 2.3850 0.1275 2.4450 0.1875 ;
        RECT 2.3850 0.8400 2.4450 0.9000 ;
        RECT 2.2800 0.4800 2.3400 0.5400 ;
        RECT 2.1750 0.2250 2.2350 0.2850 ;
        RECT 2.1750 0.7200 2.2350 0.7800 ;
        RECT 2.0700 0.4875 2.1300 0.5475 ;
        RECT 1.9650 0.1275 2.0250 0.1875 ;
        RECT 1.9650 0.8475 2.0250 0.9075 ;
        RECT 1.8600 0.4875 1.9200 0.5475 ;
        RECT 1.7550 0.2250 1.8150 0.2850 ;
        RECT 1.7550 0.7200 1.8150 0.7800 ;
        RECT 1.6500 0.4875 1.7100 0.5475 ;
        RECT 1.5450 0.1575 1.6050 0.2175 ;
        RECT 1.5450 0.6975 1.6050 0.7575 ;
        RECT 1.5450 0.8625 1.6050 0.9225 ;
        RECT 1.4400 0.4725 1.5000 0.5325 ;
        RECT 1.3350 0.7950 1.3950 0.8550 ;
        RECT 1.2300 0.4725 1.2900 0.5325 ;
        RECT 1.1250 0.1725 1.1850 0.2325 ;
        RECT 1.1250 0.8325 1.1850 0.8925 ;
        RECT 0.9150 0.1575 0.9750 0.2175 ;
        RECT 0.9150 0.8325 0.9750 0.8925 ;
        RECT 0.8175 0.4725 0.8775 0.5325 ;
        RECT 0.7050 0.6825 0.7650 0.7425 ;
        RECT 0.6000 0.4725 0.6600 0.5325 ;
        RECT 0.4950 0.1875 0.5550 0.2475 ;
        RECT 0.4950 0.8325 0.5550 0.8925 ;
        RECT 0.3900 0.4800 0.4500 0.5400 ;
        RECT 0.2850 0.6825 0.3450 0.7425 ;
        RECT 0.1800 0.4800 0.2400 0.5400 ;
        RECT 0.0750 0.1575 0.1350 0.2175 ;
        RECT 0.0750 0.8175 0.1350 0.8775 ;
        LAYER M1 ;
        RECT 2.6175 0.1500 2.6925 0.7575 ;
        RECT 2.5725 0.1500 2.6175 0.2550 ;
        RECT 2.3925 0.6825 2.6175 0.7575 ;
        RECT 2.4675 0.3300 2.5425 0.5775 ;
        RECT 2.4525 0.3300 2.4675 0.4050 ;
        RECT 2.3325 0.2625 2.4525 0.4050 ;
        RECT 2.3175 0.4800 2.3925 0.7575 ;
        RECT 1.6200 0.4800 2.3175 0.5550 ;
        RECT 2.1525 0.1950 2.2575 0.3825 ;
        RECT 2.1675 0.6300 2.2425 0.8325 ;
        RECT 1.8225 0.6300 2.1675 0.7200 ;
        RECT 1.8375 0.2925 2.1525 0.3825 ;
        RECT 1.7325 0.1950 1.8375 0.3825 ;
        RECT 1.7475 0.6300 1.8225 0.8325 ;
        RECT 1.3650 0.3225 1.5000 0.5700 ;
        RECT 1.3050 0.6525 1.4100 0.9000 ;
        RECT 0.7950 0.6525 1.3050 0.7275 ;
        RECT 1.0575 0.1500 1.2900 0.2925 ;
        RECT 1.0875 0.3675 1.2900 0.5775 ;
        RECT 0.8175 0.3900 1.0125 0.5775 ;
        RECT 0.1575 0.8250 1.0050 0.9000 ;
        RECT 0.4950 0.1500 0.8325 0.2850 ;
        RECT 0.6750 0.6525 0.7950 0.7500 ;
        RECT 0.5325 0.3825 0.7350 0.5775 ;
        RECT 0.4500 0.6750 0.5550 0.7500 ;
        RECT 0.4200 0.4425 0.4500 0.5700 ;
        RECT 0.2250 0.6450 0.4500 0.7500 ;
        RECT 0.3150 0.1500 0.4200 0.5700 ;
        RECT 0.0525 0.7950 0.1575 0.9000 ;
        LAYER VIA1 ;
        RECT 2.4675 0.4200 2.5425 0.4950 ;
        RECT 1.1325 0.1575 1.2075 0.2325 ;
        RECT 0.7125 0.1725 0.7875 0.2475 ;
        RECT 0.4275 0.6750 0.5025 0.7500 ;
        LAYER M2 ;
        RECT 2.3775 0.4200 2.5875 0.4950 ;
        RECT 2.3025 0.1125 2.3775 0.4950 ;
        RECT 1.2525 0.1125 2.3025 0.1875 ;
        RECT 1.0875 0.1125 1.2525 0.2325 ;
        RECT 0.7875 0.1125 1.0875 0.1875 ;
        RECT 0.7125 0.1125 0.7875 0.3375 ;
        RECT 0.5700 0.2625 0.7125 0.3375 ;
        RECT 0.4950 0.2625 0.5700 0.7500 ;
        RECT 0.3825 0.6750 0.4950 0.7500 ;
    END
END AOI222_0111


MACRO AOI222_1000
    CLASS CORE ;
    FOREIGN AOI222_1000 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.6800 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 0.8625 0.1125 1.0125 0.2550 ;
        RECT 0.5775 0.1125 0.8625 0.1875 ;
        RECT 0.4275 0.1125 0.5775 0.2550 ;
        RECT 0.0600 0.1125 0.4275 0.1875 ;
        VIA 0.9375 0.2025 VIA12_square ;
        VIA 0.5025 0.2025 VIA12_square ;
        END
    END ZN
    PIN C2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.5225 0.3675 1.6275 0.6375 ;
        RECT 1.4475 0.4650 1.5225 0.6375 ;
        END
    END C2
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.1325 0.2625 1.5975 0.3375 ;
        VIA 1.3350 0.3000 VIA12_square ;
        END
    END C1
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.7725 0.4125 0.8475 0.9375 ;
        RECT 0.3075 0.8625 0.7725 0.9375 ;
        VIA 0.8100 0.4950 VIA12_square ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.1400 0.8625 1.6050 0.9375 ;
        RECT 1.0650 0.4950 1.1400 0.9375 ;
        RECT 0.9750 0.4950 1.0650 0.6000 ;
        VIA 1.0575 0.5475 VIA12_square ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1425 0.3675 0.2325 0.5775 ;
        RECT 0.0675 0.3675 0.1425 0.6825 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.4575 0.7125 0.6375 0.7875 ;
        RECT 0.3825 0.4350 0.4575 0.7875 ;
        RECT 0.0675 0.7125 0.3825 0.7875 ;
        VIA 0.4200 0.5175 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.6125 -0.0750 1.6800 0.0750 ;
        RECT 1.5075 -0.0750 1.6125 0.2475 ;
        RECT 0.7875 -0.0750 1.5075 0.0750 ;
        RECT 0.6825 -0.0750 0.7875 0.2475 ;
        RECT 0.1425 -0.0750 0.6825 0.0750 ;
        RECT 0.0675 -0.0750 0.1425 0.2475 ;
        RECT 0.0000 -0.0750 0.0675 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.4250 0.9750 1.6800 1.1250 ;
        RECT 1.3050 0.8625 1.4250 1.1250 ;
        RECT 0.0000 0.9750 1.3050 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.5450 0.1575 1.6050 0.2175 ;
        RECT 1.5450 0.8175 1.6050 0.8775 ;
        RECT 1.4475 0.4950 1.5075 0.5550 ;
        RECT 1.3350 0.8700 1.3950 0.9300 ;
        RECT 1.2375 0.4725 1.2975 0.5325 ;
        RECT 1.1250 0.1725 1.1850 0.2325 ;
        RECT 1.1250 0.7800 1.1850 0.8400 ;
        RECT 1.0200 0.4725 1.0800 0.5325 ;
        RECT 0.9150 0.8325 0.9750 0.8925 ;
        RECT 0.8100 0.4725 0.8700 0.5325 ;
        RECT 0.7050 0.1575 0.7650 0.2175 ;
        RECT 0.7050 0.6675 0.7650 0.7275 ;
        RECT 0.4950 0.1575 0.5550 0.2175 ;
        RECT 0.4950 0.8325 0.5550 0.8925 ;
        RECT 0.3900 0.4800 0.4500 0.5400 ;
        RECT 0.2850 0.6825 0.3450 0.7425 ;
        RECT 0.1725 0.4800 0.2325 0.5400 ;
        RECT 0.0750 0.1575 0.1350 0.2175 ;
        RECT 0.0750 0.8175 0.1350 0.8775 ;
        LAYER M1 ;
        RECT 1.5225 0.7125 1.6275 0.9000 ;
        RECT 1.1925 0.7125 1.5225 0.7875 ;
        RECT 1.3725 0.2175 1.4025 0.3825 ;
        RECT 1.2900 0.2175 1.3725 0.5775 ;
        RECT 1.2375 0.4275 1.2900 0.5775 ;
        RECT 0.8625 0.1500 1.2150 0.2775 ;
        RECT 1.1175 0.6750 1.1925 0.8700 ;
        RECT 0.9750 0.3675 1.1625 0.6000 ;
        RECT 0.7875 0.6750 1.1175 0.7500 ;
        RECT 0.1575 0.8250 1.0050 0.9000 ;
        RECT 0.6825 0.3675 0.9000 0.5700 ;
        RECT 0.6825 0.6450 0.7875 0.7500 ;
        RECT 0.5325 0.1500 0.6075 0.7500 ;
        RECT 0.4200 0.1500 0.5325 0.2625 ;
        RECT 0.2550 0.6750 0.5325 0.7500 ;
        RECT 0.3075 0.3375 0.4575 0.6000 ;
        RECT 0.0525 0.7950 0.1575 0.9000 ;
    END
END AOI222_1000


MACRO AOI222_1010
    CLASS CORE ;
    FOREIGN AOI222_1010 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.6800 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 0.8625 0.1125 1.0125 0.2550 ;
        RECT 0.5775 0.1125 0.8625 0.1875 ;
        RECT 0.4275 0.1125 0.5775 0.2550 ;
        RECT 0.0600 0.1125 0.4275 0.1875 ;
        VIA 0.9375 0.2025 VIA12_square ;
        VIA 0.5025 0.2025 VIA12_square ;
        END
    END ZN
    PIN C2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.5225 0.3675 1.6275 0.6375 ;
        RECT 1.4475 0.4650 1.5225 0.6375 ;
        END
    END C2
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.1325 0.2625 1.5975 0.3375 ;
        VIA 1.3350 0.3000 VIA12_square ;
        END
    END C1
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.7725 0.4125 0.8475 0.9375 ;
        RECT 0.3075 0.8625 0.7725 0.9375 ;
        VIA 0.8100 0.4950 VIA12_square ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.1400 0.8625 1.6050 0.9375 ;
        RECT 1.0650 0.4950 1.1400 0.9375 ;
        RECT 0.9750 0.4950 1.0650 0.6000 ;
        VIA 1.0575 0.5475 VIA12_square ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1425 0.3675 0.2325 0.5775 ;
        RECT 0.0675 0.3675 0.1425 0.6825 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.4575 0.7125 0.6375 0.7875 ;
        RECT 0.3825 0.4350 0.4575 0.7875 ;
        RECT 0.0675 0.7125 0.3825 0.7875 ;
        VIA 0.4200 0.5175 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.6125 -0.0750 1.6800 0.0750 ;
        RECT 1.5075 -0.0750 1.6125 0.2475 ;
        RECT 0.7875 -0.0750 1.5075 0.0750 ;
        RECT 0.6825 -0.0750 0.7875 0.2475 ;
        RECT 0.1425 -0.0750 0.6825 0.0750 ;
        RECT 0.0675 -0.0750 0.1425 0.2475 ;
        RECT 0.0000 -0.0750 0.0675 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.4250 0.9750 1.6800 1.1250 ;
        RECT 1.3050 0.8625 1.4250 1.1250 ;
        RECT 0.0000 0.9750 1.3050 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.5450 0.1575 1.6050 0.2175 ;
        RECT 1.5450 0.8175 1.6050 0.8775 ;
        RECT 1.4475 0.4950 1.5075 0.5550 ;
        RECT 1.3350 0.8700 1.3950 0.9300 ;
        RECT 1.2375 0.4725 1.2975 0.5325 ;
        RECT 1.1250 0.1725 1.1850 0.2325 ;
        RECT 1.1250 0.7800 1.1850 0.8400 ;
        RECT 1.0200 0.4725 1.0800 0.5325 ;
        RECT 0.9150 0.8325 0.9750 0.8925 ;
        RECT 0.8100 0.4725 0.8700 0.5325 ;
        RECT 0.7050 0.1575 0.7650 0.2175 ;
        RECT 0.7050 0.6675 0.7650 0.7275 ;
        RECT 0.4950 0.1575 0.5550 0.2175 ;
        RECT 0.4950 0.8325 0.5550 0.8925 ;
        RECT 0.3900 0.4800 0.4500 0.5400 ;
        RECT 0.2850 0.6825 0.3450 0.7425 ;
        RECT 0.1725 0.4800 0.2325 0.5400 ;
        RECT 0.0750 0.1575 0.1350 0.2175 ;
        RECT 0.0750 0.8175 0.1350 0.8775 ;
        LAYER M1 ;
        RECT 1.5225 0.7125 1.6275 0.9000 ;
        RECT 1.1925 0.7125 1.5225 0.7875 ;
        RECT 1.3725 0.2175 1.4025 0.3825 ;
        RECT 1.2900 0.2175 1.3725 0.5775 ;
        RECT 1.2375 0.4275 1.2900 0.5775 ;
        RECT 0.8625 0.1500 1.2150 0.2775 ;
        RECT 1.1175 0.6750 1.1925 0.8700 ;
        RECT 0.9750 0.3675 1.1625 0.6000 ;
        RECT 0.7875 0.6750 1.1175 0.7500 ;
        RECT 0.1575 0.8250 1.0050 0.9000 ;
        RECT 0.6825 0.3675 0.9000 0.5700 ;
        RECT 0.6825 0.6450 0.7875 0.7500 ;
        RECT 0.5325 0.1500 0.6075 0.7500 ;
        RECT 0.4200 0.1500 0.5325 0.2625 ;
        RECT 0.2550 0.6750 0.5325 0.7500 ;
        RECT 0.3075 0.3375 0.4575 0.6000 ;
        RECT 0.0525 0.7950 0.1575 0.9000 ;
    END
END AOI222_1010


MACRO AOI22_0011
    CLASS CORE ;
    FOREIGN AOI22_0011 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.6100 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 1.1025 0.2775 3.9375 0.3975 ;
        RECT 1.1025 0.6525 1.2600 0.7725 ;
        RECT 0.7875 0.2775 1.1025 0.7725 ;
        RECT 0.6300 0.2775 0.7875 0.3975 ;
        RECT 0.6300 0.6525 0.7875 0.7725 ;
        VIA 3.7800 0.3375 VIA12_slot ;
        VIA 1.1025 0.3375 VIA12_slot ;
        VIA 1.1025 0.7125 VIA12_slot ;
        VIA 0.7875 0.3375 VIA12_slot ;
        VIA 0.7875 0.7125 VIA12_slot ;
        END
    END ZN
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 8.3100 0.4125 8.4750 0.6375 ;
        RECT 6.0375 0.4575 8.3100 0.5625 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 5.7675 0.4125 5.9325 0.6375 ;
        RECT 3.5100 0.4575 5.7675 0.5625 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 3.4050 0.5625 3.7575 0.6375 ;
        RECT 3.2700 0.4725 3.4050 0.6375 ;
        VIA 3.3375 0.5475 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1425 0.4650 1.7325 0.5550 ;
        RECT 0.0375 0.3675 0.1425 0.6825 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 8.3550 -0.0750 8.6100 0.0750 ;
        RECT 8.2350 -0.0750 8.3550 0.1875 ;
        RECT 7.9350 -0.0750 8.2350 0.0750 ;
        RECT 7.8150 -0.0750 7.9350 0.1875 ;
        RECT 7.5150 -0.0750 7.8150 0.0750 ;
        RECT 7.3950 -0.0750 7.5150 0.1875 ;
        RECT 7.0950 -0.0750 7.3950 0.0750 ;
        RECT 6.9750 -0.0750 7.0950 0.1875 ;
        RECT 6.6750 -0.0750 6.9750 0.0750 ;
        RECT 6.5550 -0.0750 6.6750 0.1875 ;
        RECT 6.2550 -0.0750 6.5550 0.0750 ;
        RECT 6.1350 -0.0750 6.2550 0.1875 ;
        RECT 3.3150 -0.0750 6.1350 0.0750 ;
        RECT 3.1950 -0.0750 3.3150 0.2250 ;
        RECT 2.8950 -0.0750 3.1950 0.0750 ;
        RECT 2.7750 -0.0750 2.8950 0.2250 ;
        RECT 2.4750 -0.0750 2.7750 0.0750 ;
        RECT 2.3550 -0.0750 2.4750 0.2250 ;
        RECT 2.0550 -0.0750 2.3550 0.0750 ;
        RECT 1.9350 -0.0750 2.0550 0.2250 ;
        RECT 0.0000 -0.0750 1.9350 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 8.3550 0.9750 8.6100 1.1250 ;
        RECT 8.2350 0.8625 8.3550 1.1250 ;
        RECT 7.9350 0.9750 8.2350 1.1250 ;
        RECT 7.8150 0.8625 7.9350 1.1250 ;
        RECT 7.5150 0.9750 7.8150 1.1250 ;
        RECT 7.3950 0.8625 7.5150 1.1250 ;
        RECT 7.0950 0.9750 7.3950 1.1250 ;
        RECT 6.9750 0.8625 7.0950 1.1250 ;
        RECT 6.6750 0.9750 6.9750 1.1250 ;
        RECT 6.5550 0.8625 6.6750 1.1250 ;
        RECT 6.2550 0.9750 6.5550 1.1250 ;
        RECT 6.1350 0.8625 6.2550 1.1250 ;
        RECT 5.8350 0.9750 6.1350 1.1250 ;
        RECT 5.7150 0.8625 5.8350 1.1250 ;
        RECT 5.4150 0.9750 5.7150 1.1250 ;
        RECT 5.2950 0.8625 5.4150 1.1250 ;
        RECT 4.9950 0.9750 5.2950 1.1250 ;
        RECT 4.8750 0.8625 4.9950 1.1250 ;
        RECT 4.5750 0.9750 4.8750 1.1250 ;
        RECT 4.4550 0.8625 4.5750 1.1250 ;
        RECT 4.1550 0.9750 4.4550 1.1250 ;
        RECT 4.0350 0.8625 4.1550 1.1250 ;
        RECT 3.7500 0.9750 4.0350 1.1250 ;
        RECT 3.6150 0.8625 3.7500 1.1250 ;
        RECT 0.0000 0.9750 3.6150 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 8.4750 0.2325 8.5350 0.2925 ;
        RECT 8.4750 0.7575 8.5350 0.8175 ;
        RECT 8.3700 0.4800 8.4300 0.5400 ;
        RECT 8.2650 0.1275 8.3250 0.1875 ;
        RECT 8.2650 0.8625 8.3250 0.9225 ;
        RECT 8.1600 0.4800 8.2200 0.5400 ;
        RECT 8.0550 0.2700 8.1150 0.3300 ;
        RECT 8.0550 0.7200 8.1150 0.7800 ;
        RECT 7.9500 0.4800 8.0100 0.5400 ;
        RECT 7.8450 0.1275 7.9050 0.1875 ;
        RECT 7.8450 0.8625 7.9050 0.9225 ;
        RECT 7.7400 0.4800 7.8000 0.5400 ;
        RECT 7.6350 0.2700 7.6950 0.3300 ;
        RECT 7.6350 0.7200 7.6950 0.7800 ;
        RECT 7.5300 0.4800 7.5900 0.5400 ;
        RECT 7.4250 0.1275 7.4850 0.1875 ;
        RECT 7.4250 0.8625 7.4850 0.9225 ;
        RECT 7.3200 0.4800 7.3800 0.5400 ;
        RECT 7.2150 0.2700 7.2750 0.3300 ;
        RECT 7.2150 0.7200 7.2750 0.7800 ;
        RECT 7.1100 0.4800 7.1700 0.5400 ;
        RECT 7.0050 0.1275 7.0650 0.1875 ;
        RECT 7.0050 0.8625 7.0650 0.9225 ;
        RECT 6.9000 0.4800 6.9600 0.5400 ;
        RECT 6.7950 0.2700 6.8550 0.3300 ;
        RECT 6.7950 0.7200 6.8550 0.7800 ;
        RECT 6.6900 0.4800 6.7500 0.5400 ;
        RECT 6.5850 0.1275 6.6450 0.1875 ;
        RECT 6.5850 0.8625 6.6450 0.9225 ;
        RECT 6.4800 0.4800 6.5400 0.5400 ;
        RECT 6.3750 0.2700 6.4350 0.3300 ;
        RECT 6.3750 0.7200 6.4350 0.7800 ;
        RECT 6.2700 0.4800 6.3300 0.5400 ;
        RECT 6.1650 0.1275 6.2250 0.1875 ;
        RECT 6.1650 0.8625 6.2250 0.9225 ;
        RECT 6.0600 0.4800 6.1200 0.5400 ;
        RECT 5.9550 0.2175 6.0150 0.2775 ;
        RECT 5.9550 0.7200 6.0150 0.7800 ;
        RECT 5.8500 0.4800 5.9100 0.5400 ;
        RECT 5.7450 0.8625 5.8050 0.9225 ;
        RECT 5.6400 0.4800 5.7000 0.5400 ;
        RECT 5.5350 0.1575 5.5950 0.2175 ;
        RECT 5.5350 0.7200 5.5950 0.7800 ;
        RECT 5.4300 0.4800 5.4900 0.5400 ;
        RECT 5.3250 0.3000 5.3850 0.3600 ;
        RECT 5.3250 0.8625 5.3850 0.9225 ;
        RECT 5.2200 0.4800 5.2800 0.5400 ;
        RECT 5.1150 0.1575 5.1750 0.2175 ;
        RECT 5.1150 0.7200 5.1750 0.7800 ;
        RECT 5.0100 0.4800 5.0700 0.5400 ;
        RECT 4.9050 0.3000 4.9650 0.3600 ;
        RECT 4.9050 0.8625 4.9650 0.9225 ;
        RECT 4.8000 0.4800 4.8600 0.5400 ;
        RECT 4.6950 0.1575 4.7550 0.2175 ;
        RECT 4.6950 0.7200 4.7550 0.7800 ;
        RECT 4.5900 0.4800 4.6500 0.5400 ;
        RECT 4.4850 0.3000 4.5450 0.3600 ;
        RECT 4.4850 0.8625 4.5450 0.9225 ;
        RECT 4.3800 0.4800 4.4400 0.5400 ;
        RECT 4.2750 0.1575 4.3350 0.2175 ;
        RECT 4.2750 0.7200 4.3350 0.7800 ;
        RECT 4.1700 0.4800 4.2300 0.5400 ;
        RECT 4.0650 0.3000 4.1250 0.3600 ;
        RECT 4.0650 0.8625 4.1250 0.9225 ;
        RECT 3.9600 0.4800 4.0200 0.5400 ;
        RECT 3.8550 0.1575 3.9150 0.2175 ;
        RECT 3.8550 0.7200 3.9150 0.7800 ;
        RECT 3.7500 0.4800 3.8100 0.5400 ;
        RECT 3.6450 0.8625 3.7050 0.9225 ;
        RECT 3.5400 0.4875 3.6000 0.5475 ;
        RECT 3.4350 0.2325 3.4950 0.2925 ;
        RECT 3.4350 0.7800 3.4950 0.8400 ;
        RECT 3.3300 0.4800 3.3900 0.5400 ;
        RECT 3.2250 0.1500 3.2850 0.2100 ;
        RECT 3.2250 0.6825 3.2850 0.7425 ;
        RECT 3.1200 0.4800 3.1800 0.5400 ;
        RECT 3.0150 0.2325 3.0750 0.2925 ;
        RECT 3.0150 0.8325 3.0750 0.8925 ;
        RECT 2.9100 0.4800 2.9700 0.5400 ;
        RECT 2.8050 0.1500 2.8650 0.2100 ;
        RECT 2.8050 0.6825 2.8650 0.7425 ;
        RECT 2.7000 0.4800 2.7600 0.5400 ;
        RECT 2.5950 0.2325 2.6550 0.2925 ;
        RECT 2.5950 0.8325 2.6550 0.8925 ;
        RECT 2.4900 0.4800 2.5500 0.5400 ;
        RECT 2.3850 0.1500 2.4450 0.2100 ;
        RECT 2.3850 0.6825 2.4450 0.7425 ;
        RECT 2.2800 0.4800 2.3400 0.5400 ;
        RECT 2.1750 0.2325 2.2350 0.2925 ;
        RECT 2.1750 0.8325 2.2350 0.8925 ;
        RECT 2.0700 0.4800 2.1300 0.5400 ;
        RECT 1.9650 0.1500 2.0250 0.2100 ;
        RECT 1.9650 0.6825 2.0250 0.7425 ;
        RECT 1.8675 0.4800 1.9275 0.5400 ;
        RECT 1.7550 0.2250 1.8150 0.2850 ;
        RECT 1.7550 0.8325 1.8150 0.8925 ;
        RECT 1.6425 0.4875 1.7025 0.5475 ;
        RECT 1.5450 0.3075 1.6050 0.3675 ;
        RECT 1.5450 0.6825 1.6050 0.7425 ;
        RECT 1.4400 0.4875 1.5000 0.5475 ;
        RECT 1.3350 0.1575 1.3950 0.2175 ;
        RECT 1.3350 0.8250 1.3950 0.8850 ;
        RECT 1.2300 0.4875 1.2900 0.5475 ;
        RECT 1.1250 0.3075 1.1850 0.3675 ;
        RECT 1.1250 0.6825 1.1850 0.7425 ;
        RECT 1.0200 0.4875 1.0800 0.5475 ;
        RECT 0.9150 0.1575 0.9750 0.2175 ;
        RECT 0.9150 0.8250 0.9750 0.8850 ;
        RECT 0.8100 0.4875 0.8700 0.5475 ;
        RECT 0.7050 0.3075 0.7650 0.3675 ;
        RECT 0.7050 0.6825 0.7650 0.7425 ;
        RECT 0.6000 0.4800 0.6600 0.5400 ;
        RECT 0.4950 0.1575 0.5550 0.2175 ;
        RECT 0.4950 0.8250 0.5550 0.8850 ;
        RECT 0.3900 0.4800 0.4500 0.5400 ;
        RECT 0.2850 0.3075 0.3450 0.3675 ;
        RECT 0.2850 0.6675 0.3450 0.7275 ;
        RECT 0.1800 0.4800 0.2400 0.5400 ;
        RECT 0.0750 0.1725 0.1350 0.2325 ;
        RECT 0.0750 0.8175 0.1350 0.8775 ;
        LAYER M1 ;
        RECT 8.4675 0.1875 8.5425 0.3375 ;
        RECT 8.4675 0.7125 8.5425 0.8625 ;
        RECT 6.0225 0.2625 8.4675 0.3375 ;
        RECT 3.5025 0.7125 8.4675 0.7875 ;
        RECT 5.9475 0.1500 6.0225 0.3375 ;
        RECT 3.8175 0.1500 5.9475 0.2250 ;
        RECT 3.6075 0.3000 5.4300 0.3750 ;
        RECT 3.4275 0.1875 3.5025 0.3750 ;
        RECT 3.4275 0.7125 3.5025 0.9000 ;
        RECT 3.0825 0.3000 3.4275 0.3750 ;
        RECT 0.1575 0.8250 3.4275 0.9000 ;
        RECT 3.2550 0.4725 3.4200 0.6000 ;
        RECT 0.3825 0.6750 3.3150 0.7500 ;
        RECT 1.8375 0.4725 3.2550 0.5475 ;
        RECT 3.0075 0.1875 3.0825 0.3750 ;
        RECT 2.6625 0.3000 3.0075 0.3750 ;
        RECT 2.5875 0.1875 2.6625 0.3750 ;
        RECT 2.2425 0.3000 2.5875 0.3750 ;
        RECT 2.1675 0.1875 2.2425 0.3750 ;
        RECT 1.8225 0.3000 2.1675 0.3750 ;
        RECT 1.7475 0.1500 1.8225 0.3750 ;
        RECT 0.1575 0.1500 1.7475 0.2250 ;
        RECT 0.2550 0.3000 1.6425 0.3900 ;
        RECT 0.2625 0.6450 0.3825 0.7500 ;
        RECT 0.0525 0.1500 0.1575 0.2550 ;
        RECT 0.0525 0.7950 0.1575 0.9000 ;
        LAYER M2 ;
        RECT 1.1325 0.2775 3.9375 0.3975 ;
        RECT 1.1325 0.6525 1.2600 0.7725 ;
        RECT 0.6300 0.2775 0.7575 0.3975 ;
        RECT 0.6300 0.6525 0.7575 0.7725 ;
    END
END AOI22_0011


MACRO AOI22_0111
    CLASS CORE ;
    FOREIGN AOI22_0111 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.7800 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 0.6825 0.2850 2.4600 0.3900 ;
        RECT 0.3675 0.2850 0.6825 0.7800 ;
        VIA 2.3025 0.3375 VIA12_slot ;
        VIA 0.5250 0.3450 VIA12_slot ;
        VIA 0.5250 0.7125 VIA12_slot ;
        END
    END ZN
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 2.8875 0.5625 3.3525 0.6375 ;
        VIA 3.1275 0.6000 VIA12_square ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 2.1975 0.5625 2.6625 0.6375 ;
        VIA 2.4150 0.6000 VIA12_square ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.5825 0.5625 2.0475 0.6375 ;
        VIA 1.8300 0.6000 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1425 0.4650 0.8925 0.5550 ;
        RECT 0.0375 0.3675 0.1425 0.6825 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 3.5250 -0.0750 3.7800 0.0750 ;
        RECT 3.4050 -0.0750 3.5250 0.1875 ;
        RECT 3.1050 -0.0750 3.4050 0.0750 ;
        RECT 2.9850 -0.0750 3.1050 0.1875 ;
        RECT 1.6350 -0.0750 2.9850 0.0750 ;
        RECT 1.5150 -0.0750 1.6350 0.2250 ;
        RECT 1.2150 -0.0750 1.5150 0.0750 ;
        RECT 1.0950 -0.0750 1.2150 0.2250 ;
        RECT 0.0000 -0.0750 1.0950 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 3.5250 0.9750 3.7800 1.1250 ;
        RECT 3.4050 0.8625 3.5250 1.1250 ;
        RECT 3.1050 0.9750 3.4050 1.1250 ;
        RECT 2.9850 0.8625 3.1050 1.1250 ;
        RECT 2.6850 0.9750 2.9850 1.1250 ;
        RECT 2.5650 0.8625 2.6850 1.1250 ;
        RECT 2.2650 0.9750 2.5650 1.1250 ;
        RECT 2.1450 0.8625 2.2650 1.1250 ;
        RECT 0.0000 0.9750 2.1450 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 3.6450 0.2475 3.7050 0.3075 ;
        RECT 3.6450 0.7500 3.7050 0.8100 ;
        RECT 3.5400 0.4800 3.6000 0.5400 ;
        RECT 3.4350 0.1275 3.4950 0.1875 ;
        RECT 3.4350 0.8700 3.4950 0.9300 ;
        RECT 3.3300 0.4800 3.3900 0.5400 ;
        RECT 3.2250 0.2700 3.2850 0.3300 ;
        RECT 3.2250 0.7200 3.2850 0.7800 ;
        RECT 3.1200 0.4800 3.1800 0.5400 ;
        RECT 3.0150 0.1275 3.0750 0.1875 ;
        RECT 3.0150 0.8700 3.0750 0.9300 ;
        RECT 2.9100 0.4800 2.9700 0.5400 ;
        RECT 2.8050 0.2175 2.8650 0.2775 ;
        RECT 2.8050 0.7200 2.8650 0.7800 ;
        RECT 2.7000 0.4800 2.7600 0.5400 ;
        RECT 2.5950 0.3000 2.6550 0.3600 ;
        RECT 2.5950 0.8700 2.6550 0.9300 ;
        RECT 2.4900 0.4800 2.5500 0.5400 ;
        RECT 2.3850 0.1575 2.4450 0.2175 ;
        RECT 2.3850 0.7200 2.4450 0.7800 ;
        RECT 2.2800 0.4800 2.3400 0.5400 ;
        RECT 2.1750 0.3000 2.2350 0.3600 ;
        RECT 2.1750 0.8700 2.2350 0.9300 ;
        RECT 2.0700 0.4800 2.1300 0.5400 ;
        RECT 1.9650 0.1575 2.0250 0.2175 ;
        RECT 1.9650 0.7200 2.0250 0.7800 ;
        RECT 1.7550 0.3000 1.8150 0.3600 ;
        RECT 1.7550 0.8325 1.8150 0.8925 ;
        RECT 1.6500 0.4800 1.7100 0.5400 ;
        RECT 1.5450 0.1500 1.6050 0.2100 ;
        RECT 1.5450 0.6825 1.6050 0.7425 ;
        RECT 1.4400 0.4800 1.5000 0.5400 ;
        RECT 1.3350 0.3000 1.3950 0.3600 ;
        RECT 1.3350 0.8325 1.3950 0.8925 ;
        RECT 1.2300 0.4800 1.2900 0.5400 ;
        RECT 1.1250 0.1500 1.1850 0.2100 ;
        RECT 1.1250 0.6825 1.1850 0.7425 ;
        RECT 1.0275 0.4800 1.0875 0.5400 ;
        RECT 0.9150 0.2250 0.9750 0.2850 ;
        RECT 0.9150 0.8325 0.9750 0.8925 ;
        RECT 0.8025 0.4875 0.8625 0.5475 ;
        RECT 0.7050 0.3075 0.7650 0.3675 ;
        RECT 0.7050 0.6825 0.7650 0.7425 ;
        RECT 0.6000 0.4800 0.6600 0.5400 ;
        RECT 0.4950 0.1575 0.5550 0.2175 ;
        RECT 0.4950 0.8250 0.5550 0.8850 ;
        RECT 0.3900 0.4800 0.4500 0.5400 ;
        RECT 0.2850 0.3075 0.3450 0.3675 ;
        RECT 0.2850 0.6675 0.3450 0.7275 ;
        RECT 0.1800 0.4800 0.2400 0.5400 ;
        RECT 0.0750 0.1800 0.1350 0.2400 ;
        RECT 0.0750 0.8175 0.1350 0.8775 ;
        LAYER M1 ;
        RECT 3.6375 0.2175 3.7125 0.3375 ;
        RECT 3.6225 0.7125 3.7125 0.8475 ;
        RECT 2.8725 0.2625 3.6375 0.3375 ;
        RECT 3.2100 0.4575 3.6375 0.5625 ;
        RECT 1.8600 0.7125 3.6225 0.7875 ;
        RECT 3.0450 0.4575 3.2100 0.6375 ;
        RECT 2.8875 0.4575 3.0450 0.5625 ;
        RECT 2.7975 0.1500 2.8725 0.3375 ;
        RECT 1.9350 0.1500 2.7975 0.2250 ;
        RECT 2.4975 0.4575 2.7825 0.5625 ;
        RECT 2.0700 0.3000 2.6925 0.3750 ;
        RECT 2.3325 0.4575 2.4975 0.6375 ;
        RECT 2.0475 0.4575 2.3325 0.5625 ;
        RECT 1.7475 0.4725 1.9125 0.6375 ;
        RECT 1.7700 0.7125 1.8600 0.9000 ;
        RECT 0.9825 0.3000 1.8450 0.3750 ;
        RECT 0.1575 0.8250 1.7700 0.9000 ;
        RECT 0.9975 0.4725 1.7475 0.5475 ;
        RECT 0.3825 0.6750 1.6350 0.7500 ;
        RECT 0.9075 0.1500 0.9825 0.3750 ;
        RECT 0.1425 0.1500 0.9075 0.2250 ;
        RECT 0.2475 0.3000 0.8025 0.3900 ;
        RECT 0.2625 0.6450 0.3825 0.7500 ;
        RECT 0.0525 0.7950 0.1575 0.9000 ;
        RECT 0.0375 0.1500 0.1425 0.2700 ;
        LAYER M2 ;
        RECT 0.7125 0.2850 2.4600 0.3900 ;
    END
END AOI22_0111


MACRO AOI22_1000
    CLASS CORE ;
    FOREIGN AOI22_1000 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.0500 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 0.4650 0.8625 0.8700 0.9375 ;
        RECT 0.3600 0.5700 0.4650 0.9375 ;
        VIA 0.4125 0.6450 VIA12_square ;
        END
    END ZN
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.9075 0.3675 1.0125 0.6375 ;
        RECT 0.8175 0.4725 0.9075 0.6375 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.4800 0.2625 0.9450 0.3375 ;
        VIA 0.7050 0.3000 VIA12_square ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.1500 0.4125 0.6225 0.4875 ;
        VIA 0.2625 0.4500 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.3600 0.1125 0.7200 0.1875 ;
        RECT 0.2550 0.1125 0.3600 0.2775 ;
        VIA 0.3075 0.1950 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.0050 -0.0750 1.0500 0.0750 ;
        RECT 0.8850 -0.0750 1.0050 0.2925 ;
        RECT 0.1200 -0.0750 0.8850 0.0750 ;
        RECT 0.1200 0.2700 0.1500 0.3975 ;
        RECT 0.0450 -0.0750 0.1200 0.3975 ;
        RECT 0.0000 -0.0750 0.0450 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.7950 0.9750 1.0500 1.1250 ;
        RECT 0.6750 0.8625 0.7950 1.1250 ;
        RECT 0.0000 0.9750 0.6750 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 0.9150 0.2325 0.9750 0.2925 ;
        RECT 0.9150 0.8175 0.9750 0.8775 ;
        RECT 0.8175 0.5025 0.8775 0.5625 ;
        RECT 0.7050 0.8700 0.7650 0.9300 ;
        RECT 0.6000 0.5100 0.6600 0.5700 ;
        RECT 0.4950 0.3300 0.5550 0.3900 ;
        RECT 0.4950 0.8325 0.5550 0.8925 ;
        RECT 0.3900 0.1500 0.4500 0.2100 ;
        RECT 0.2850 0.6825 0.3450 0.7425 ;
        RECT 0.1800 0.4875 0.2400 0.5475 ;
        RECT 0.0750 0.3075 0.1350 0.3675 ;
        RECT 0.0750 0.8250 0.1350 0.8850 ;
        LAYER M1 ;
        RECT 0.8925 0.7125 0.9975 0.9000 ;
        RECT 0.6000 0.7125 0.8925 0.7875 ;
        RECT 0.6675 0.1800 0.7425 0.6150 ;
        RECT 0.5625 0.5100 0.6675 0.6150 ;
        RECT 0.5250 0.7125 0.6000 0.9000 ;
        RECT 0.4500 0.3300 0.5925 0.4350 ;
        RECT 0.2250 0.1500 0.5550 0.2550 ;
        RECT 0.1425 0.8250 0.5250 0.9000 ;
        RECT 0.3750 0.3300 0.4500 0.7500 ;
        RECT 0.2550 0.6450 0.3750 0.7500 ;
        RECT 0.2250 0.3600 0.3000 0.5700 ;
        RECT 0.1650 0.4725 0.2250 0.5700 ;
        RECT 0.0600 0.4725 0.1650 0.6450 ;
        RECT 0.0375 0.7950 0.1425 0.9000 ;
    END
END AOI22_1000


MACRO AOI22_1010
    CLASS CORE ;
    FOREIGN AOI22_1010 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.0500 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.4500 0.3300 0.5925 0.4350 ;
        RECT 0.3750 0.3300 0.4500 0.7500 ;
        RECT 0.2625 0.6450 0.3750 0.7500 ;
        END
    END ZN
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.9075 0.3675 1.0125 0.6375 ;
        RECT 0.8175 0.4725 0.9075 0.6375 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.6675 0.1800 0.7425 0.6375 ;
        RECT 0.5625 0.5100 0.6675 0.6375 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.2250 0.3600 0.3000 0.5700 ;
        RECT 0.1650 0.4725 0.2250 0.5700 ;
        RECT 0.0600 0.4725 0.1650 0.6825 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.3600 0.1125 0.5925 0.1875 ;
        RECT 0.2550 0.1125 0.3600 0.2775 ;
        RECT 0.1275 0.1125 0.2550 0.1875 ;
        VIA 0.3075 0.1950 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.0050 -0.0750 1.0500 0.0750 ;
        RECT 0.8850 -0.0750 1.0050 0.2625 ;
        RECT 0.1200 -0.0750 0.8850 0.0750 ;
        RECT 0.1200 0.2700 0.1500 0.3975 ;
        RECT 0.0450 -0.0750 0.1200 0.3975 ;
        RECT 0.0000 -0.0750 0.0450 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.7950 0.9750 1.0500 1.1250 ;
        RECT 0.6750 0.8625 0.7950 1.1250 ;
        RECT 0.0000 0.9750 0.6750 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 0.9150 0.1875 0.9750 0.2475 ;
        RECT 0.9150 0.7725 0.9750 0.8325 ;
        RECT 0.8175 0.5025 0.8775 0.5625 ;
        RECT 0.7050 0.8700 0.7650 0.9300 ;
        RECT 0.6000 0.5100 0.6600 0.5700 ;
        RECT 0.4950 0.3300 0.5550 0.3900 ;
        RECT 0.4950 0.8325 0.5550 0.8925 ;
        RECT 0.3900 0.1500 0.4500 0.2100 ;
        RECT 0.2850 0.6675 0.3450 0.7275 ;
        RECT 0.1800 0.4875 0.2400 0.5475 ;
        RECT 0.0750 0.3075 0.1350 0.3675 ;
        RECT 0.0750 0.8250 0.1350 0.8850 ;
        LAYER M1 ;
        RECT 0.8925 0.7125 0.9825 0.8700 ;
        RECT 0.6000 0.7125 0.8925 0.7875 ;
        RECT 0.5250 0.7125 0.6000 0.9000 ;
        RECT 0.2250 0.1500 0.5550 0.2550 ;
        RECT 0.1425 0.8250 0.5250 0.9000 ;
        RECT 0.0375 0.7950 0.1425 0.9000 ;
    END
END AOI22_1010


MACRO AOI31_0011
    CLASS CORE ;
    FOREIGN AOI31_0011 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.8900 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 1.4850 0.1125 1.6350 0.2550 ;
        RECT 1.2225 0.1125 1.4850 0.1875 ;
        RECT 1.1475 0.1125 1.2225 0.7875 ;
        RECT 0.6825 0.7125 1.1475 0.7875 ;
        VIA 1.5600 0.2025 VIA12_square ;
        VIA 1.1850 0.2250 VIA12_square ;
        VIA 1.1850 0.6975 VIA12_square ;
        END
    END ZN
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.7475 0.3675 1.8225 0.6375 ;
        RECT 1.6575 0.4500 1.7475 0.6375 ;
        RECT 1.4475 0.4500 1.6575 0.5700 ;
        END
    END B
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.2975 0.3975 1.3725 0.9375 ;
        RECT 0.4275 0.8625 1.2975 0.9375 ;
        RECT 0.3525 0.4125 0.4275 0.9375 ;
        RECT 0.1425 0.4125 0.3525 0.4875 ;
        VIA 1.3350 0.4875 VIA12_square ;
        VIA 0.2250 0.4500 VIA12_square ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.3825 0.2625 0.8475 0.3375 ;
        VIA 0.4950 0.3000 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.8100 0.5625 1.0275 0.6375 ;
        RECT 0.6600 0.4650 0.8100 0.6375 ;
        RECT 0.5475 0.5625 0.6600 0.6375 ;
        VIA 0.7350 0.5175 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.8225 -0.0750 1.8900 0.0750 ;
        RECT 1.7475 -0.0750 1.8225 0.2625 ;
        RECT 1.4025 -0.0750 1.7475 0.0750 ;
        RECT 1.3275 -0.0750 1.4025 0.2700 ;
        RECT 0.1575 -0.0750 1.3275 0.0750 ;
        RECT 0.0525 -0.0750 0.1575 0.3000 ;
        RECT 0.0000 -0.0750 0.0525 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.6350 0.9750 1.8900 1.1250 ;
        RECT 1.5150 0.8625 1.6350 1.1250 ;
        RECT 0.0000 0.9750 1.5150 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.7550 0.1725 1.8150 0.2325 ;
        RECT 1.7550 0.7350 1.8150 0.7950 ;
        RECT 1.6500 0.4800 1.7100 0.5400 ;
        RECT 1.5450 0.2325 1.6050 0.2925 ;
        RECT 1.5450 0.8700 1.6050 0.9300 ;
        RECT 1.4475 0.4800 1.5075 0.5400 ;
        RECT 1.3350 0.1800 1.3950 0.2400 ;
        RECT 1.3350 0.8325 1.3950 0.8925 ;
        RECT 1.2300 0.4800 1.2900 0.5400 ;
        RECT 1.1250 0.6675 1.1850 0.7275 ;
        RECT 1.0200 0.4800 1.0800 0.5400 ;
        RECT 0.9150 0.8325 0.9750 0.8925 ;
        RECT 0.8100 0.4875 0.8700 0.5475 ;
        RECT 0.7050 0.1650 0.7650 0.2250 ;
        RECT 0.7050 0.6675 0.7650 0.7275 ;
        RECT 0.6000 0.4875 0.6600 0.5475 ;
        RECT 0.4950 0.8325 0.5550 0.8925 ;
        RECT 0.3900 0.4800 0.4500 0.5400 ;
        RECT 0.2850 0.6675 0.3450 0.7275 ;
        RECT 0.1800 0.4725 0.2400 0.5325 ;
        RECT 0.0750 0.2100 0.1350 0.2700 ;
        RECT 0.0750 0.8175 0.1350 0.8775 ;
        LAYER M1 ;
        RECT 1.7325 0.7125 1.8375 0.8175 ;
        RECT 1.4400 0.7125 1.7325 0.7875 ;
        RECT 1.4775 0.1500 1.6725 0.3150 ;
        RECT 1.3650 0.7125 1.4400 0.9000 ;
        RECT 1.1625 0.3750 1.3725 0.5700 ;
        RECT 0.1575 0.8250 1.3650 0.9000 ;
        RECT 0.2550 0.6450 1.2675 0.7500 ;
        RECT 1.1325 0.1500 1.2375 0.3000 ;
        RECT 0.6750 0.1500 1.1325 0.2400 ;
        RECT 1.0425 0.4500 1.0875 0.5700 ;
        RECT 0.9675 0.3150 1.0425 0.5700 ;
        RECT 0.5625 0.3150 0.9675 0.3900 ;
        RECT 0.5775 0.4650 0.8925 0.5700 ;
        RECT 0.5025 0.2175 0.5625 0.3900 ;
        RECT 0.4275 0.2175 0.5025 0.5700 ;
        RECT 0.3825 0.4500 0.4275 0.5700 ;
        RECT 0.1050 0.3750 0.3075 0.5700 ;
        RECT 0.0525 0.7950 0.1575 0.9000 ;
    END
END AOI31_0011


MACRO AOI31_0111
    CLASS CORE ;
    FOREIGN AOI31_0111 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.7800 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 0.3675 0.2850 0.6825 0.7575 ;
        VIA 0.5250 0.3450 VIA12_slot ;
        VIA 0.5250 0.6975 VIA12_slot ;
        END
    END ZN
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 3.6375 0.3675 3.7125 0.6375 ;
        RECT 3.5475 0.4650 3.6375 0.6375 ;
        RECT 2.9025 0.4650 3.5475 0.5850 ;
        END
    END B
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 2.2425 0.4125 2.5575 0.4875 ;
        RECT 2.1675 0.4125 2.2425 0.6375 ;
        RECT 1.8525 0.5625 2.1675 0.6375 ;
        VIA 2.2050 0.5175 VIA12_square ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.4025 0.5625 1.7175 0.6375 ;
        RECT 1.3275 0.4125 1.4025 0.6375 ;
        RECT 1.0125 0.4125 1.3275 0.4875 ;
        VIA 1.3650 0.5175 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1425 0.4650 0.8925 0.5700 ;
        RECT 0.0675 0.3675 0.1425 0.6825 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 3.7125 -0.0750 3.7800 0.0750 ;
        RECT 3.6375 -0.0750 3.7125 0.2625 ;
        RECT 3.3150 -0.0750 3.6375 0.0750 ;
        RECT 3.1950 -0.0750 3.3150 0.2100 ;
        RECT 2.8950 -0.0750 3.1950 0.0750 ;
        RECT 2.7750 -0.0750 2.8950 0.2100 ;
        RECT 2.4675 -0.0750 2.7750 0.0750 ;
        RECT 2.3625 -0.0750 2.4675 0.2400 ;
        RECT 2.0550 -0.0750 2.3625 0.0750 ;
        RECT 1.9500 -0.0750 2.0550 0.2475 ;
        RECT 0.0000 -0.0750 1.9500 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 3.5250 0.9750 3.7800 1.1250 ;
        RECT 3.4050 0.8625 3.5250 1.1250 ;
        RECT 3.0975 0.9750 3.4050 1.1250 ;
        RECT 2.9925 0.8100 3.0975 1.1250 ;
        RECT 0.0000 0.9750 2.9925 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 3.6450 0.1725 3.7050 0.2325 ;
        RECT 3.6450 0.7350 3.7050 0.7950 ;
        RECT 3.5400 0.4950 3.6000 0.5550 ;
        RECT 3.4350 0.3075 3.4950 0.3675 ;
        RECT 3.4350 0.8700 3.4950 0.9300 ;
        RECT 3.3300 0.4950 3.3900 0.5550 ;
        RECT 3.2250 0.1425 3.2850 0.2025 ;
        RECT 3.2250 0.6975 3.2850 0.7575 ;
        RECT 3.1200 0.4950 3.1800 0.5550 ;
        RECT 3.0150 0.3075 3.0750 0.3675 ;
        RECT 3.0150 0.8325 3.0750 0.8925 ;
        RECT 2.9100 0.4950 2.9700 0.5550 ;
        RECT 2.8050 0.1425 2.8650 0.2025 ;
        RECT 2.8050 0.7425 2.8650 0.8025 ;
        RECT 2.7000 0.4950 2.7600 0.5550 ;
        RECT 2.5950 0.2475 2.6550 0.3075 ;
        RECT 2.5950 0.6675 2.6550 0.7275 ;
        RECT 2.4900 0.4950 2.5500 0.5550 ;
        RECT 2.3850 0.1575 2.4450 0.2175 ;
        RECT 2.3850 0.8325 2.4450 0.8925 ;
        RECT 2.2800 0.4950 2.3400 0.5550 ;
        RECT 2.1750 0.3225 2.2350 0.3825 ;
        RECT 2.1750 0.6675 2.2350 0.7275 ;
        RECT 2.0700 0.4950 2.1300 0.5550 ;
        RECT 1.9650 0.1575 2.0250 0.2175 ;
        RECT 1.9650 0.8325 2.0250 0.8925 ;
        RECT 1.7550 0.1575 1.8150 0.2175 ;
        RECT 1.7550 0.8325 1.8150 0.8925 ;
        RECT 1.6500 0.4875 1.7100 0.5475 ;
        RECT 1.5450 0.3150 1.6050 0.3750 ;
        RECT 1.5450 0.6675 1.6050 0.7275 ;
        RECT 1.4400 0.4875 1.5000 0.5475 ;
        RECT 1.3350 0.1575 1.3950 0.2175 ;
        RECT 1.3350 0.8325 1.3950 0.8925 ;
        RECT 1.2300 0.4875 1.2900 0.5475 ;
        RECT 1.1250 0.3150 1.1850 0.3750 ;
        RECT 1.1250 0.6675 1.1850 0.7275 ;
        RECT 1.0200 0.4875 1.0800 0.5475 ;
        RECT 0.9150 0.1575 0.9750 0.2175 ;
        RECT 0.9150 0.8325 0.9750 0.8925 ;
        RECT 0.8100 0.4875 0.8700 0.5475 ;
        RECT 0.7050 0.3150 0.7650 0.3750 ;
        RECT 0.7050 0.6675 0.7650 0.7275 ;
        RECT 0.6000 0.4875 0.6600 0.5475 ;
        RECT 0.4950 0.1575 0.5550 0.2175 ;
        RECT 0.4950 0.8325 0.5550 0.8925 ;
        RECT 0.3900 0.4875 0.4500 0.5475 ;
        RECT 0.2850 0.3150 0.3450 0.3750 ;
        RECT 0.2850 0.6675 0.3450 0.7275 ;
        RECT 0.1800 0.4875 0.2400 0.5475 ;
        RECT 0.0750 0.1800 0.1350 0.2400 ;
        RECT 0.0750 0.8175 0.1350 0.8775 ;
        LAYER M1 ;
        RECT 3.6225 0.7125 3.7275 0.8175 ;
        RECT 3.3225 0.7125 3.6225 0.7875 ;
        RECT 2.7525 0.2850 3.5175 0.3900 ;
        RECT 3.1875 0.6600 3.3225 0.7875 ;
        RECT 2.8725 0.6600 3.1875 0.7350 ;
        RECT 2.7975 0.6600 2.8725 0.9000 ;
        RECT 0.1575 0.8250 2.7975 0.9000 ;
        RECT 2.0400 0.4725 2.7900 0.5700 ;
        RECT 0.2550 0.6450 2.7225 0.7500 ;
        RECT 2.5875 0.2100 2.6625 0.3975 ;
        RECT 1.8900 0.3225 2.5875 0.3975 ;
        RECT 1.8150 0.3075 1.8900 0.3975 ;
        RECT 0.1575 0.1500 1.8450 0.2250 ;
        RECT 1.0950 0.3075 1.8150 0.3825 ;
        RECT 0.9975 0.4650 1.7325 0.5700 ;
        RECT 0.2550 0.3000 0.7950 0.3900 ;
        RECT 0.0525 0.1500 0.1575 0.2625 ;
        RECT 0.0525 0.7950 0.1575 0.9000 ;
        LAYER VIA1 ;
        RECT 2.8425 0.3000 2.9175 0.3750 ;
        RECT 2.6025 0.6600 2.6775 0.7350 ;
        LAYER M2 ;
        RECT 2.8725 0.3000 2.9925 0.3750 ;
        RECT 2.7975 0.3000 2.8725 0.7500 ;
        RECT 2.5575 0.6450 2.7975 0.7500 ;
    END
END AOI31_0111


MACRO AOI31_1000
    CLASS CORE ;
    FOREIGN AOI31_1000 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.2600 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.9450 0.1500 1.0050 0.3825 ;
        RECT 0.8700 0.1500 0.9450 0.7425 ;
        RECT 0.6750 0.1500 0.8700 0.2550 ;
        RECT 0.2550 0.6675 0.8700 0.7425 ;
        END
    END ZN
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.1175 0.3675 1.1925 0.6825 ;
        RECT 1.0200 0.4800 1.1175 0.6000 ;
        END
    END B
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1425 0.4500 0.2400 0.5700 ;
        RECT 0.0675 0.3675 0.1425 0.6825 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.3900 0.4500 0.4500 0.5700 ;
        RECT 0.3150 0.2175 0.3900 0.5700 ;
        RECT 0.2775 0.2175 0.3150 0.3825 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.6000 0.3675 0.7725 0.5325 ;
        RECT 0.5250 0.2175 0.6000 0.5325 ;
        RECT 0.4875 0.2175 0.5250 0.3825 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.2075 -0.0750 1.2600 0.0750 ;
        RECT 1.1025 -0.0750 1.2075 0.2475 ;
        RECT 0.1650 -0.0750 1.1025 0.0750 ;
        RECT 0.0450 -0.0750 0.1650 0.2325 ;
        RECT 0.0000 -0.0750 0.0450 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.2150 0.9750 1.2600 1.1250 ;
        RECT 1.1100 0.8025 1.2150 1.1250 ;
        RECT 0.0000 0.9750 1.1100 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.1250 0.1575 1.1850 0.2175 ;
        RECT 1.1250 0.8325 1.1850 0.8925 ;
        RECT 1.0200 0.5100 1.0800 0.5700 ;
        RECT 0.9150 0.1575 0.9750 0.2175 ;
        RECT 0.9150 0.8325 0.9750 0.8925 ;
        RECT 0.7050 0.1575 0.7650 0.2175 ;
        RECT 0.7050 0.6750 0.7650 0.7350 ;
        RECT 0.6000 0.4650 0.6600 0.5250 ;
        RECT 0.4950 0.8325 0.5550 0.8925 ;
        RECT 0.3900 0.4800 0.4500 0.5400 ;
        RECT 0.2850 0.6750 0.3450 0.7350 ;
        RECT 0.1800 0.4800 0.2400 0.5400 ;
        RECT 0.0750 0.1575 0.1350 0.2175 ;
        RECT 0.0750 0.8175 0.1350 0.8775 ;
        LAYER M1 ;
        RECT 0.1575 0.8250 1.0050 0.9000 ;
        RECT 0.0525 0.7950 0.1575 0.9000 ;
    END
END AOI31_1000


MACRO AOI31_1010
    CLASS CORE ;
    FOREIGN AOI31_1010 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.2600 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.9450 0.1500 0.9825 0.3825 ;
        RECT 0.8700 0.1500 0.9450 0.7425 ;
        RECT 0.7050 0.1500 0.8700 0.2700 ;
        RECT 0.2550 0.6675 0.8700 0.7425 ;
        END
    END ZN
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.1175 0.3675 1.1925 0.6825 ;
        RECT 1.0200 0.4575 1.1175 0.5775 ;
        END
    END B
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1425 0.4500 0.2400 0.5700 ;
        RECT 0.0675 0.3675 0.1425 0.6825 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.3900 0.4500 0.4500 0.5700 ;
        RECT 0.3150 0.2175 0.3900 0.5700 ;
        RECT 0.2775 0.2175 0.3150 0.3825 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.6000 0.3675 0.7725 0.5325 ;
        RECT 0.5250 0.2175 0.6000 0.5325 ;
        RECT 0.4875 0.2175 0.5250 0.3825 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.2075 -0.0750 1.2600 0.0750 ;
        RECT 1.1025 -0.0750 1.2075 0.2625 ;
        RECT 0.1650 -0.0750 1.1025 0.0750 ;
        RECT 0.0450 -0.0750 0.1650 0.2325 ;
        RECT 0.0000 -0.0750 0.0450 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.2150 0.9750 1.2600 1.1250 ;
        RECT 1.1100 0.8025 1.2150 1.1250 ;
        RECT 0.0000 0.9750 1.1100 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.1250 0.1725 1.1850 0.2325 ;
        RECT 1.1250 0.8325 1.1850 0.8925 ;
        RECT 1.0200 0.4875 1.0800 0.5475 ;
        RECT 0.9150 0.2325 0.9750 0.2925 ;
        RECT 0.9150 0.8325 0.9750 0.8925 ;
        RECT 0.7050 0.1800 0.7650 0.2400 ;
        RECT 0.7050 0.6750 0.7650 0.7350 ;
        RECT 0.6000 0.4650 0.6600 0.5250 ;
        RECT 0.4950 0.8325 0.5550 0.8925 ;
        RECT 0.3900 0.4800 0.4500 0.5400 ;
        RECT 0.2850 0.6750 0.3450 0.7350 ;
        RECT 0.1800 0.4800 0.2400 0.5400 ;
        RECT 0.0750 0.1575 0.1350 0.2175 ;
        RECT 0.0750 0.8175 0.1350 0.8775 ;
        LAYER M1 ;
        RECT 0.1575 0.8250 1.0050 0.9000 ;
        RECT 0.0525 0.7950 0.1575 0.9000 ;
    END
END AOI31_1010


MACRO AOI32_0011
    CLASS CORE ;
    FOREIGN AOI32_0011 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.3100 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 1.5150 0.1125 1.6650 0.2550 ;
        RECT 1.2225 0.1125 1.5150 0.1875 ;
        RECT 1.1475 0.1125 1.2225 0.7875 ;
        RECT 0.6825 0.7125 1.1475 0.7875 ;
        VIA 1.5900 0.2025 VIA12_square ;
        VIA 1.1850 0.2250 VIA12_square ;
        VIA 1.1850 0.6975 VIA12_square ;
        END
    END ZN
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 2.0625 0.3150 2.2425 0.6375 ;
        RECT 1.5525 0.3150 2.0625 0.3900 ;
        RECT 1.4700 0.3150 1.5525 0.5700 ;
        RECT 1.4475 0.4500 1.4700 0.5700 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.7850 0.8625 2.2500 0.9375 ;
        RECT 1.7100 0.4425 1.7850 0.9375 ;
        RECT 1.6800 0.4425 1.7100 0.5925 ;
        VIA 1.7325 0.5175 VIA12_square ;
        END
    END B1
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.2975 0.4050 1.3725 0.9375 ;
        RECT 0.4275 0.8625 1.2975 0.9375 ;
        RECT 0.3525 0.4125 0.4275 0.9375 ;
        RECT 0.1425 0.4125 0.3525 0.4875 ;
        VIA 1.3350 0.4875 VIA12_square ;
        VIA 0.2550 0.4500 VIA12_square ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.3900 0.2625 0.8550 0.3375 ;
        VIA 0.5025 0.3000 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.8100 0.5625 1.0275 0.6375 ;
        RECT 0.6600 0.4650 0.8100 0.6375 ;
        RECT 0.5475 0.5625 0.6600 0.6375 ;
        VIA 0.7350 0.5175 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 2.2650 -0.0750 2.3100 0.0750 ;
        RECT 2.1450 -0.0750 2.2650 0.2250 ;
        RECT 1.4025 -0.0750 2.1450 0.0750 ;
        RECT 1.3275 -0.0750 1.4025 0.2625 ;
        RECT 0.1575 -0.0750 1.3275 0.0750 ;
        RECT 0.0525 -0.0750 0.1575 0.2925 ;
        RECT 0.0000 -0.0750 0.0525 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 2.0550 0.9750 2.3100 1.1250 ;
        RECT 1.9350 0.8625 2.0550 1.1250 ;
        RECT 1.6275 0.9750 1.9350 1.1250 ;
        RECT 1.5225 0.8025 1.6275 1.1250 ;
        RECT 0.0000 0.9750 1.5225 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 2.1750 0.1575 2.2350 0.2175 ;
        RECT 2.1750 0.7350 2.2350 0.7950 ;
        RECT 2.0700 0.4800 2.1300 0.5400 ;
        RECT 1.9650 0.8700 2.0250 0.9300 ;
        RECT 1.8600 0.4875 1.9200 0.5475 ;
        RECT 1.7550 0.1650 1.8150 0.2250 ;
        RECT 1.7550 0.6900 1.8150 0.7500 ;
        RECT 1.6500 0.4875 1.7100 0.5475 ;
        RECT 1.5450 0.8250 1.6050 0.8850 ;
        RECT 1.4475 0.4800 1.5075 0.5400 ;
        RECT 1.3350 0.1725 1.3950 0.2325 ;
        RECT 1.3350 0.8325 1.3950 0.8925 ;
        RECT 1.2300 0.4800 1.2900 0.5400 ;
        RECT 1.1250 0.6675 1.1850 0.7275 ;
        RECT 1.0200 0.4800 1.0800 0.5400 ;
        RECT 0.9150 0.8325 0.9750 0.8925 ;
        RECT 0.8100 0.4875 0.8700 0.5475 ;
        RECT 0.7050 0.1650 0.7650 0.2250 ;
        RECT 0.7050 0.6675 0.7650 0.7275 ;
        RECT 0.6000 0.4875 0.6600 0.5475 ;
        RECT 0.4950 0.8325 0.5550 0.8925 ;
        RECT 0.3900 0.4800 0.4500 0.5400 ;
        RECT 0.2850 0.6675 0.3450 0.7275 ;
        RECT 0.1800 0.4725 0.2400 0.5325 ;
        RECT 0.0750 0.2100 0.1350 0.2700 ;
        RECT 0.0750 0.8175 0.1350 0.8775 ;
        LAYER M1 ;
        RECT 2.1525 0.7125 2.2575 0.8175 ;
        RECT 1.8300 0.7125 2.1525 0.7875 ;
        RECT 1.6275 0.4650 1.9425 0.5700 ;
        RECT 1.5075 0.1500 1.8675 0.2400 ;
        RECT 1.7400 0.6525 1.8300 0.7875 ;
        RECT 1.4475 0.6525 1.7400 0.7275 ;
        RECT 1.3725 0.6525 1.4475 0.9000 ;
        RECT 1.1625 0.3750 1.3725 0.5700 ;
        RECT 0.1575 0.8250 1.3725 0.9000 ;
        RECT 0.2550 0.6450 1.2600 0.7500 ;
        RECT 1.1325 0.1500 1.2375 0.3000 ;
        RECT 0.6750 0.1500 1.1325 0.2400 ;
        RECT 1.0575 0.4500 1.0875 0.5700 ;
        RECT 0.9825 0.3150 1.0575 0.5700 ;
        RECT 0.5625 0.3150 0.9825 0.3900 ;
        RECT 0.5775 0.4650 0.8925 0.5700 ;
        RECT 0.5025 0.2175 0.5625 0.3900 ;
        RECT 0.4275 0.2175 0.5025 0.5700 ;
        RECT 0.3825 0.4500 0.4275 0.5700 ;
        RECT 0.1125 0.3675 0.3075 0.5700 ;
        RECT 0.0525 0.7950 0.1575 0.9000 ;
    END
END AOI32_0011


MACRO AOI32_0111
    CLASS CORE ;
    FOREIGN AOI32_0111 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.5200 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 1.6275 0.2625 1.9425 0.7650 ;
        VIA 1.7850 0.3450 VIA12_slot ;
        VIA 1.7850 0.6825 VIA12_slot ;
        END
    END ZN
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.3125 0.8625 1.7025 0.9375 ;
        RECT 1.2375 0.4725 1.3125 0.9375 ;
        VIA 1.2750 0.5550 VIA12_square ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.9975 0.2625 1.4625 0.3375 ;
        VIA 1.0875 0.3000 VIA12_square ;
        END
    END B1
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.1125 0.4125 0.5775 0.4875 ;
        VIA 0.2400 0.4500 VIA12_square ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.1125 0.2625 0.5775 0.3375 ;
        VIA 0.4200 0.3000 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.9225 0.4125 0.9525 0.5775 ;
        RECT 0.8475 0.4125 0.9225 0.9375 ;
        RECT 0.3825 0.8625 0.8475 0.9375 ;
        VIA 0.9000 0.4950 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 2.2650 -0.0750 2.5200 0.0750 ;
        RECT 2.1450 -0.0750 2.2650 0.1875 ;
        RECT 1.8450 -0.0750 2.1450 0.0750 ;
        RECT 1.7250 -0.0750 1.8450 0.1950 ;
        RECT 1.4175 -0.0750 1.7250 0.0750 ;
        RECT 1.3125 -0.0750 1.4175 0.2325 ;
        RECT 0.1425 -0.0750 1.3125 0.0750 ;
        RECT 0.0675 -0.0750 0.1425 0.2550 ;
        RECT 0.0000 -0.0750 0.0675 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 2.2650 0.9750 2.5200 1.1250 ;
        RECT 2.1450 0.8325 2.2650 1.1250 ;
        RECT 1.8225 0.9750 2.1450 1.1250 ;
        RECT 1.7475 0.8250 1.8225 1.1250 ;
        RECT 1.4175 0.9750 1.7475 1.1250 ;
        RECT 1.3125 0.8100 1.4175 1.1250 ;
        RECT 1.0050 0.9750 1.3125 1.1250 ;
        RECT 0.8850 0.8325 1.0050 1.1250 ;
        RECT 0.0000 0.9750 0.8850 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 2.3850 0.1725 2.4450 0.2325 ;
        RECT 2.3850 0.6900 2.4450 0.7500 ;
        RECT 2.2725 0.4650 2.3325 0.5250 ;
        RECT 2.1750 0.1275 2.2350 0.1875 ;
        RECT 2.1750 0.8400 2.2350 0.9000 ;
        RECT 2.0700 0.4800 2.1300 0.5400 ;
        RECT 1.9650 0.2250 2.0250 0.2850 ;
        RECT 1.9650 0.7200 2.0250 0.7800 ;
        RECT 1.8600 0.4800 1.9200 0.5400 ;
        RECT 1.7550 0.1275 1.8150 0.1875 ;
        RECT 1.7550 0.8550 1.8150 0.9150 ;
        RECT 1.6500 0.4800 1.7100 0.5400 ;
        RECT 1.5450 0.2250 1.6050 0.2850 ;
        RECT 1.5450 0.7200 1.6050 0.7800 ;
        RECT 1.4400 0.4800 1.5000 0.5400 ;
        RECT 1.3350 0.1425 1.3950 0.2025 ;
        RECT 1.3350 0.8325 1.3950 0.8925 ;
        RECT 1.2300 0.4950 1.2900 0.5550 ;
        RECT 1.1250 0.7800 1.1850 0.8400 ;
        RECT 1.0275 0.4725 1.0875 0.5325 ;
        RECT 0.9150 0.1800 0.9750 0.2400 ;
        RECT 0.9150 0.8325 0.9750 0.8925 ;
        RECT 0.7050 0.2025 0.7650 0.2625 ;
        RECT 0.7050 0.8325 0.7650 0.8925 ;
        RECT 0.6000 0.4800 0.6600 0.5400 ;
        RECT 0.4950 0.6825 0.5550 0.7425 ;
        RECT 0.3900 0.4950 0.4500 0.5550 ;
        RECT 0.2850 0.8325 0.3450 0.8925 ;
        RECT 0.1800 0.4950 0.2400 0.5550 ;
        RECT 0.0750 0.1575 0.1350 0.2175 ;
        RECT 0.0750 0.7575 0.1350 0.8175 ;
        LAYER M1 ;
        RECT 2.4075 0.1500 2.4825 0.7575 ;
        RECT 2.3625 0.1500 2.4075 0.2550 ;
        RECT 2.1825 0.6825 2.4075 0.7575 ;
        RECT 2.2575 0.3300 2.3325 0.5775 ;
        RECT 2.2425 0.3300 2.2575 0.4050 ;
        RECT 2.1075 0.2625 2.2425 0.4050 ;
        RECT 2.1075 0.4800 2.1825 0.7575 ;
        RECT 1.5225 0.4800 2.1075 0.5625 ;
        RECT 1.9425 0.1950 2.0325 0.3825 ;
        RECT 1.9575 0.6375 2.0325 0.8325 ;
        RECT 1.6125 0.6375 1.9575 0.7200 ;
        RECT 1.6275 0.2925 1.9425 0.3825 ;
        RECT 1.5225 0.1950 1.6275 0.3825 ;
        RECT 1.5375 0.6375 1.6125 0.8325 ;
        RECT 1.4100 0.4575 1.5225 0.5625 ;
        RECT 1.2225 0.3075 1.3350 0.6375 ;
        RECT 1.1550 0.7575 1.2075 0.8625 ;
        RECT 1.0800 0.6825 1.1550 0.8625 ;
        RECT 1.0500 0.1800 1.1400 0.5775 ;
        RECT 0.8025 0.6825 1.0800 0.7575 ;
        RECT 1.0275 0.3300 1.0500 0.5775 ;
        RECT 0.8625 0.1500 0.9750 0.2700 ;
        RECT 0.8475 0.4125 0.9525 0.5775 ;
        RECT 0.6600 0.1500 0.8625 0.3375 ;
        RECT 0.5775 0.4575 0.8475 0.5775 ;
        RECT 0.7275 0.6825 0.8025 0.9000 ;
        RECT 0.2550 0.8250 0.7275 0.9000 ;
        RECT 0.1425 0.6750 0.5850 0.7500 ;
        RECT 0.3675 0.2175 0.4725 0.5775 ;
        RECT 0.2175 0.2100 0.2925 0.6000 ;
        RECT 0.1800 0.3675 0.2175 0.6000 ;
        RECT 0.0675 0.6750 0.1425 0.8475 ;
        LAYER VIA1 ;
        RECT 2.2575 0.4200 2.3325 0.4950 ;
        RECT 0.6975 0.1950 0.7725 0.2700 ;
        RECT 0.4650 0.6750 0.5400 0.7500 ;
        LAYER M2 ;
        RECT 2.1675 0.4200 2.3775 0.4950 ;
        RECT 2.0925 0.1125 2.1675 0.4950 ;
        RECT 0.7725 0.1125 2.0925 0.1875 ;
        RECT 0.6975 0.1125 0.7725 0.7500 ;
        RECT 0.4200 0.6750 0.6975 0.7500 ;
    END
END AOI32_0111


MACRO AOI32_1000
    CLASS CORE ;
    FOREIGN AOI32_1000 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.4700 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 0.7725 0.2625 0.8925 0.3375 ;
        RECT 0.6975 0.2625 0.7725 0.9375 ;
        RECT 0.2325 0.8625 0.6975 0.9375 ;
        VIA 0.7800 0.3000 VIA12_square ;
        VIA 0.7350 0.7125 VIA12_square ;
        END
    END ZN
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.3125 0.3675 1.4175 0.6375 ;
        RECT 1.1850 0.4875 1.3125 0.6375 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.0725 0.1125 1.1775 0.3075 ;
        RECT 0.6075 0.1125 1.0725 0.1875 ;
        VIA 1.1250 0.2325 VIA12_square ;
        END
    END B1
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.1125 0.4125 0.5775 0.4875 ;
        VIA 0.2400 0.4500 VIA12_square ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.1125 0.2625 0.5775 0.3375 ;
        VIA 0.4200 0.3000 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.9225 0.8625 1.3875 0.9375 ;
        RECT 0.9225 0.4125 0.9525 0.5775 ;
        RECT 0.8475 0.4125 0.9225 0.9375 ;
        VIA 0.9000 0.4950 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.4175 -0.0750 1.4700 0.0750 ;
        RECT 1.3125 -0.0750 1.4175 0.2475 ;
        RECT 0.1425 -0.0750 1.3125 0.0750 ;
        RECT 0.0675 -0.0750 0.1425 0.2550 ;
        RECT 0.0000 -0.0750 0.0675 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.2150 0.9750 1.4700 1.1250 ;
        RECT 1.0950 0.8625 1.2150 1.1250 ;
        RECT 0.0000 0.9750 1.0950 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.3350 0.1575 1.3950 0.2175 ;
        RECT 1.3350 0.8175 1.3950 0.8775 ;
        RECT 1.2300 0.4950 1.2900 0.5550 ;
        RECT 1.1250 0.8625 1.1850 0.9225 ;
        RECT 1.0275 0.4725 1.0875 0.5325 ;
        RECT 0.9150 0.1575 0.9750 0.2175 ;
        RECT 0.9150 0.8325 0.9750 0.8925 ;
        RECT 0.7050 0.1575 0.7650 0.2175 ;
        RECT 0.7050 0.8325 0.7650 0.8925 ;
        RECT 0.6000 0.4800 0.6600 0.5400 ;
        RECT 0.4950 0.6900 0.5550 0.7500 ;
        RECT 0.3900 0.4950 0.4500 0.5550 ;
        RECT 0.2850 0.8325 0.3450 0.8925 ;
        RECT 0.1800 0.4950 0.2400 0.5550 ;
        RECT 0.0750 0.1575 0.1350 0.2175 ;
        RECT 0.0750 0.7800 0.1350 0.8400 ;
        LAYER M1 ;
        RECT 1.3125 0.7125 1.4175 0.9000 ;
        RECT 1.0200 0.7125 1.3125 0.7875 ;
        RECT 1.1100 0.1500 1.1850 0.4050 ;
        RECT 1.0800 0.1500 1.1100 0.5625 ;
        RECT 1.0275 0.3300 1.0800 0.5625 ;
        RECT 0.9450 0.7125 1.0200 0.9000 ;
        RECT 0.8625 0.1500 1.0050 0.2550 ;
        RECT 0.8475 0.4125 0.9525 0.5775 ;
        RECT 0.2550 0.8250 0.9450 0.9000 ;
        RECT 0.6600 0.1500 0.8625 0.3375 ;
        RECT 0.5775 0.4575 0.8475 0.5775 ;
        RECT 0.1425 0.6750 0.8175 0.7500 ;
        RECT 0.3675 0.2175 0.4725 0.5775 ;
        RECT 0.2175 0.2100 0.2925 0.6000 ;
        RECT 0.1800 0.3675 0.2175 0.6000 ;
        RECT 0.0675 0.6750 0.1425 0.8700 ;
    END
END AOI32_1000


MACRO AOI32_1010
    CLASS CORE ;
    FOREIGN AOI32_1010 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.4700 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 0.7725 0.2625 0.8925 0.3375 ;
        RECT 0.6975 0.2625 0.7725 0.9375 ;
        RECT 0.2325 0.8625 0.6975 0.9375 ;
        VIA 0.7800 0.3000 VIA12_square ;
        VIA 0.7350 0.7125 VIA12_square ;
        END
    END ZN
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.3125 0.3675 1.4175 0.6375 ;
        RECT 1.1850 0.4875 1.3125 0.6375 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.0725 0.1125 1.1775 0.3075 ;
        RECT 0.6075 0.1125 1.0725 0.1875 ;
        VIA 1.1250 0.2325 VIA12_square ;
        END
    END B1
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.1125 0.4125 0.5775 0.4875 ;
        VIA 0.2400 0.4500 VIA12_square ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.1125 0.2625 0.5775 0.3375 ;
        VIA 0.4200 0.3000 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.9225 0.8625 1.3875 0.9375 ;
        RECT 0.9225 0.4125 0.9525 0.5775 ;
        RECT 0.8475 0.4125 0.9225 0.9375 ;
        VIA 0.9000 0.4950 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.4175 -0.0750 1.4700 0.0750 ;
        RECT 1.3125 -0.0750 1.4175 0.2775 ;
        RECT 0.1425 -0.0750 1.3125 0.0750 ;
        RECT 0.0675 -0.0750 0.1425 0.2550 ;
        RECT 0.0000 -0.0750 0.0675 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.2150 0.9750 1.4700 1.1250 ;
        RECT 1.0950 0.8625 1.2150 1.1250 ;
        RECT 0.0000 0.9750 1.0950 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.3350 0.1875 1.3950 0.2475 ;
        RECT 1.3350 0.7425 1.3950 0.8025 ;
        RECT 1.2300 0.4950 1.2900 0.5550 ;
        RECT 1.1250 0.8625 1.1850 0.9225 ;
        RECT 1.0275 0.4725 1.0875 0.5325 ;
        RECT 0.9150 0.1725 0.9750 0.2325 ;
        RECT 0.9150 0.8325 0.9750 0.8925 ;
        RECT 0.7050 0.2025 0.7650 0.2625 ;
        RECT 0.7050 0.8325 0.7650 0.8925 ;
        RECT 0.6000 0.4800 0.6600 0.5400 ;
        RECT 0.4950 0.6825 0.5550 0.7425 ;
        RECT 0.3900 0.4950 0.4500 0.5550 ;
        RECT 0.2850 0.8325 0.3450 0.8925 ;
        RECT 0.1800 0.4950 0.2400 0.5550 ;
        RECT 0.0750 0.1575 0.1350 0.2175 ;
        RECT 0.0750 0.7575 0.1350 0.8175 ;
        LAYER M1 ;
        RECT 1.3200 0.7125 1.4100 0.8325 ;
        RECT 1.0200 0.7125 1.3200 0.7875 ;
        RECT 1.1100 0.1500 1.1775 0.4050 ;
        RECT 1.0725 0.1500 1.1100 0.5625 ;
        RECT 1.0275 0.3300 1.0725 0.5625 ;
        RECT 0.9450 0.7125 1.0200 0.9000 ;
        RECT 0.9450 0.1500 0.9975 0.2550 ;
        RECT 0.8475 0.4125 0.9525 0.5775 ;
        RECT 0.6600 0.1500 0.9450 0.3375 ;
        RECT 0.2550 0.8250 0.9450 0.9000 ;
        RECT 0.5775 0.4575 0.8475 0.5775 ;
        RECT 0.1425 0.6750 0.8175 0.7500 ;
        RECT 0.3675 0.2175 0.4725 0.5775 ;
        RECT 0.2175 0.2100 0.2925 0.6000 ;
        RECT 0.1800 0.3675 0.2175 0.6000 ;
        RECT 0.0675 0.6750 0.1425 0.8475 ;
    END
END AOI32_1010


MACRO AOI33_0011
    CLASS CORE ;
    FOREIGN AOI33_0011 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.7300 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 1.5225 0.1125 1.6875 0.2550 ;
        RECT 1.2075 0.1125 1.5225 0.1875 ;
        RECT 1.1325 0.1125 1.2075 0.7875 ;
        RECT 1.0125 0.1650 1.1325 0.2400 ;
        RECT 0.6675 0.7125 1.1325 0.7875 ;
        VIA 1.6050 0.2025 VIA12_square ;
        VIA 1.1700 0.6975 VIA12_square ;
        VIA 1.1250 0.2025 VIA12_square ;
        END
    END ZN
    PIN B3
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 2.3775 0.5625 2.6325 0.6375 ;
        RECT 2.3025 0.5625 2.3775 0.7875 ;
        RECT 1.6125 0.7125 2.3025 0.7875 ;
        RECT 1.5375 0.4050 1.6125 0.7875 ;
        RECT 1.4775 0.4050 1.5375 0.5700 ;
        VIA 2.5200 0.6000 VIA12_square ;
        VIA 1.5300 0.4875 VIA12_square ;
        END
    END B3
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.9125 0.2625 2.3775 0.3375 ;
        VIA 2.2350 0.3000 VIA12_square ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 2.0700 0.4125 2.3250 0.4875 ;
        RECT 1.9200 0.4125 2.0700 0.5700 ;
        RECT 1.8000 0.4125 1.9200 0.4875 ;
        VIA 1.9950 0.5175 VIA12_square ;
        END
    END B1
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.2825 0.4050 1.3575 0.9375 ;
        RECT 0.4275 0.8625 1.2825 0.9375 ;
        RECT 0.3525 0.4125 0.4275 0.9375 ;
        RECT 0.1575 0.4125 0.3525 0.4875 ;
        VIA 1.3200 0.4875 VIA12_square ;
        VIA 0.2700 0.4500 VIA12_square ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.3825 0.2625 0.8475 0.3375 ;
        VIA 0.4950 0.3000 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.8100 0.5625 1.0125 0.6375 ;
        RECT 0.6600 0.4650 0.8100 0.6375 ;
        RECT 0.5475 0.5625 0.6600 0.6375 ;
        VIA 0.7350 0.5175 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 2.6775 -0.0750 2.7300 0.0750 ;
        RECT 2.5725 -0.0750 2.6775 0.3000 ;
        RECT 1.4175 -0.0750 2.5725 0.0750 ;
        RECT 1.3125 -0.0750 1.4175 0.2700 ;
        RECT 0.1575 -0.0750 1.3125 0.0750 ;
        RECT 0.0525 -0.0750 0.1575 0.2925 ;
        RECT 0.0000 -0.0750 0.0525 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 2.4750 0.9750 2.7300 1.1250 ;
        RECT 2.3550 0.8625 2.4750 1.1250 ;
        RECT 2.0475 0.9750 2.3550 1.1250 ;
        RECT 1.9425 0.8025 2.0475 1.1250 ;
        RECT 1.6275 0.9750 1.9425 1.1250 ;
        RECT 1.5225 0.8025 1.6275 1.1250 ;
        RECT 0.0000 0.9750 1.5225 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 2.5950 0.2175 2.6550 0.2775 ;
        RECT 2.5950 0.7350 2.6550 0.7950 ;
        RECT 2.4900 0.4800 2.5500 0.5400 ;
        RECT 2.3850 0.8700 2.4450 0.9300 ;
        RECT 2.2800 0.4800 2.3400 0.5400 ;
        RECT 2.1750 0.6900 2.2350 0.7500 ;
        RECT 2.0700 0.4875 2.1300 0.5475 ;
        RECT 1.9650 0.1650 2.0250 0.2250 ;
        RECT 1.9650 0.8250 2.0250 0.8850 ;
        RECT 1.8600 0.4875 1.9200 0.5475 ;
        RECT 1.7550 0.6600 1.8150 0.7200 ;
        RECT 1.6500 0.4800 1.7100 0.5400 ;
        RECT 1.5450 0.8250 1.6050 0.8850 ;
        RECT 1.4400 0.4800 1.5000 0.5400 ;
        RECT 1.3350 0.1800 1.3950 0.2400 ;
        RECT 1.3350 0.7500 1.3950 0.8100 ;
        RECT 1.2300 0.4800 1.2900 0.5400 ;
        RECT 1.1250 0.6675 1.1850 0.7275 ;
        RECT 1.0200 0.4800 1.0800 0.5400 ;
        RECT 0.9150 0.8325 0.9750 0.8925 ;
        RECT 0.8100 0.4875 0.8700 0.5475 ;
        RECT 0.7050 0.1650 0.7650 0.2250 ;
        RECT 0.7050 0.6675 0.7650 0.7275 ;
        RECT 0.6000 0.4875 0.6600 0.5475 ;
        RECT 0.4950 0.8325 0.5550 0.8925 ;
        RECT 0.3900 0.4800 0.4500 0.5400 ;
        RECT 0.2850 0.6675 0.3450 0.7275 ;
        RECT 0.1800 0.4725 0.2400 0.5325 ;
        RECT 0.0750 0.2100 0.1350 0.2700 ;
        RECT 0.0750 0.8175 0.1350 0.8775 ;
        LAYER M1 ;
        RECT 2.5725 0.7125 2.6775 0.8175 ;
        RECT 2.4225 0.4050 2.6175 0.6375 ;
        RECT 2.2500 0.7125 2.5725 0.7875 ;
        RECT 2.3025 0.4500 2.3475 0.5700 ;
        RECT 2.2275 0.2175 2.3025 0.5700 ;
        RECT 2.1600 0.6525 2.2500 0.7875 ;
        RECT 2.1675 0.2175 2.2275 0.3900 ;
        RECT 1.7625 0.3150 2.1675 0.3900 ;
        RECT 1.4025 0.6525 2.1600 0.7275 ;
        RECT 1.8375 0.4650 2.1525 0.5700 ;
        RECT 1.5225 0.1500 2.0550 0.2400 ;
        RECT 1.6875 0.3150 1.7625 0.5700 ;
        RECT 1.6500 0.4500 1.6875 0.5700 ;
        RECT 1.4325 0.3450 1.5750 0.5775 ;
        RECT 1.3275 0.6525 1.4025 0.9000 ;
        RECT 1.1625 0.3450 1.3575 0.5700 ;
        RECT 0.1575 0.8250 1.3275 0.9000 ;
        RECT 0.2550 0.6450 1.2450 0.7500 ;
        RECT 0.6750 0.1500 1.2075 0.2400 ;
        RECT 1.0575 0.4500 1.0875 0.5700 ;
        RECT 0.9825 0.3150 1.0575 0.5700 ;
        RECT 0.5625 0.3150 0.9825 0.3900 ;
        RECT 0.5775 0.4650 0.8925 0.5700 ;
        RECT 0.5025 0.2175 0.5625 0.3900 ;
        RECT 0.4275 0.2175 0.5025 0.5700 ;
        RECT 0.3825 0.4500 0.4275 0.5700 ;
        RECT 0.1125 0.3675 0.3075 0.5700 ;
        RECT 0.0525 0.7950 0.1575 0.9000 ;
    END
END AOI33_0011


MACRO AOI33_0111
    CLASS CORE ;
    FOREIGN AOI33_0111 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.5200 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 1.6275 0.2625 1.9425 0.7575 ;
        VIA 1.7850 0.3450 VIA12_slot ;
        VIA 1.7850 0.6750 VIA12_slot ;
        END
    END ZN
    PIN B3
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.0275 0.7125 1.4925 0.7875 ;
        VIA 1.3800 0.7500 VIA12_square ;
        END
    END B3
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.0125 0.4125 1.4775 0.4875 ;
        VIA 1.1250 0.4500 VIA12_square ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.9000 0.2625 1.3500 0.3375 ;
        RECT 0.8250 0.2625 0.9000 0.3675 ;
        VIA 0.9375 0.3000 VIA12_square ;
        END
    END B1
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.0600 0.4125 0.5250 0.4875 ;
        VIA 0.2400 0.4500 VIA12_square ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.0600 0.2625 0.5250 0.3375 ;
        VIA 0.4125 0.3000 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.7500 0.5625 1.1775 0.6375 ;
        RECT 0.6450 0.4125 0.7500 0.6375 ;
        VIA 0.6975 0.4950 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 2.2650 -0.0750 2.5200 0.0750 ;
        RECT 2.1450 -0.0750 2.2650 0.1875 ;
        RECT 1.8450 -0.0750 2.1450 0.0750 ;
        RECT 1.7250 -0.0750 1.8450 0.1950 ;
        RECT 1.4175 -0.0750 1.7250 0.0750 ;
        RECT 1.3125 -0.0750 1.4175 0.2175 ;
        RECT 0.1425 -0.0750 1.3125 0.0750 ;
        RECT 0.0675 -0.0750 0.1425 0.2550 ;
        RECT 0.0000 -0.0750 0.0675 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 2.2650 0.9750 2.5200 1.1250 ;
        RECT 2.1450 0.8325 2.2650 1.1250 ;
        RECT 1.8225 0.9750 2.1450 1.1250 ;
        RECT 1.7475 0.8175 1.8225 1.1250 ;
        RECT 1.4250 0.9750 1.7475 1.1250 ;
        RECT 1.3050 0.8625 1.4250 1.1250 ;
        RECT 1.0050 0.9750 1.3050 1.1250 ;
        RECT 0.8850 0.8625 1.0050 1.1250 ;
        RECT 0.0000 0.9750 0.8850 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 2.3850 0.1725 2.4450 0.2325 ;
        RECT 2.3850 0.6900 2.4450 0.7500 ;
        RECT 2.2725 0.4650 2.3325 0.5250 ;
        RECT 2.1750 0.1275 2.2350 0.1875 ;
        RECT 2.1750 0.8400 2.2350 0.9000 ;
        RECT 2.0700 0.4800 2.1300 0.5400 ;
        RECT 1.9650 0.2250 2.0250 0.2850 ;
        RECT 1.9650 0.7200 2.0250 0.7800 ;
        RECT 1.8600 0.4800 1.9200 0.5400 ;
        RECT 1.7550 0.1275 1.8150 0.1875 ;
        RECT 1.7550 0.8475 1.8150 0.9075 ;
        RECT 1.6500 0.4800 1.7100 0.5400 ;
        RECT 1.5450 0.2250 1.6050 0.2850 ;
        RECT 1.5450 0.7200 1.6050 0.7800 ;
        RECT 1.4400 0.4800 1.5000 0.5400 ;
        RECT 1.3350 0.1275 1.3950 0.1875 ;
        RECT 1.3350 0.8700 1.3950 0.9300 ;
        RECT 1.2375 0.4800 1.2975 0.5400 ;
        RECT 1.1250 0.8175 1.1850 0.8775 ;
        RECT 1.0200 0.4950 1.0800 0.5550 ;
        RECT 0.9150 0.8625 0.9750 0.9225 ;
        RECT 0.8175 0.4725 0.8775 0.5325 ;
        RECT 0.7050 0.1725 0.7650 0.2325 ;
        RECT 0.7050 0.8325 0.7650 0.8925 ;
        RECT 0.6000 0.4800 0.6600 0.5400 ;
        RECT 0.4950 0.6825 0.5550 0.7425 ;
        RECT 0.3900 0.4950 0.4500 0.5550 ;
        RECT 0.2850 0.8325 0.3450 0.8925 ;
        RECT 0.1800 0.4950 0.2400 0.5550 ;
        RECT 0.0750 0.1575 0.1350 0.2175 ;
        RECT 0.0750 0.7575 0.1350 0.8175 ;
        LAYER M1 ;
        RECT 2.4075 0.1500 2.4825 0.7575 ;
        RECT 2.3625 0.1500 2.4075 0.2550 ;
        RECT 2.1825 0.6825 2.4075 0.7575 ;
        RECT 2.2575 0.3300 2.3325 0.5775 ;
        RECT 2.2425 0.3300 2.2575 0.4050 ;
        RECT 2.1075 0.2625 2.2425 0.4050 ;
        RECT 2.1075 0.4800 2.1825 0.7575 ;
        RECT 1.5225 0.4800 2.1075 0.5550 ;
        RECT 1.9425 0.1950 2.0325 0.3825 ;
        RECT 1.9575 0.6300 2.0325 0.8325 ;
        RECT 1.6125 0.6300 1.9575 0.7200 ;
        RECT 1.6275 0.2925 1.9425 0.3825 ;
        RECT 1.5225 0.1950 1.6275 0.3825 ;
        RECT 1.5375 0.6300 1.6125 0.8325 ;
        RECT 1.4100 0.4575 1.5225 0.5550 ;
        RECT 1.3125 0.6375 1.4625 0.7875 ;
        RECT 1.2975 0.4350 1.3125 0.7875 ;
        RECT 1.2375 0.4350 1.2975 0.7125 ;
        RECT 1.1550 0.7950 1.2075 0.9000 ;
        RECT 1.0575 0.3225 1.1625 0.5850 ;
        RECT 1.0800 0.7125 1.1550 0.9000 ;
        RECT 0.8100 0.7125 1.0800 0.7875 ;
        RECT 0.9900 0.4800 1.0575 0.5850 ;
        RECT 0.9000 0.1800 0.9825 0.4050 ;
        RECT 0.8625 0.1800 0.9000 0.5625 ;
        RECT 0.8175 0.3300 0.8625 0.5625 ;
        RECT 0.7350 0.7125 0.8100 0.9000 ;
        RECT 0.6900 0.1500 0.7875 0.2550 ;
        RECT 0.5475 0.4125 0.7425 0.6000 ;
        RECT 0.2550 0.8250 0.7350 0.9000 ;
        RECT 0.5475 0.1500 0.6900 0.3375 ;
        RECT 0.1425 0.6750 0.6225 0.7500 ;
        RECT 0.3675 0.2175 0.4725 0.5775 ;
        RECT 0.2175 0.2100 0.2925 0.6000 ;
        RECT 0.1800 0.3675 0.2175 0.6000 ;
        RECT 0.0675 0.6750 0.1425 0.8475 ;
        LAYER VIA1 ;
        RECT 2.2575 0.4200 2.3325 0.4950 ;
        RECT 0.6600 0.1650 0.7350 0.2400 ;
        RECT 0.4425 0.6750 0.5175 0.7500 ;
        LAYER M2 ;
        RECT 2.1675 0.4200 2.3775 0.4950 ;
        RECT 2.0925 0.1125 2.1675 0.9375 ;
        RECT 0.7500 0.1125 2.0925 0.1875 ;
        RECT 0.5325 0.8625 2.0925 0.9375 ;
        RECT 0.6450 0.1125 0.7500 0.2775 ;
        RECT 0.4275 0.6375 0.5325 0.9375 ;
    END
END AOI33_0111


MACRO AOI33_1000
    CLASS CORE ;
    FOREIGN AOI33_1000 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.6800 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 0.7725 0.2625 0.8625 0.3375 ;
        RECT 0.6975 0.2625 0.7725 0.9375 ;
        RECT 0.2325 0.8625 0.6975 0.9375 ;
        VIA 0.7800 0.3000 VIA12_square ;
        VIA 0.7350 0.7125 VIA12_square ;
        END
    END ZN
    PIN B3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.5225 0.3675 1.6275 0.6825 ;
        RECT 1.4475 0.4500 1.5225 0.5700 ;
        END
    END B3
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.2825 0.7125 1.6200 0.7875 ;
        RECT 1.1775 0.4725 1.2825 0.7875 ;
        RECT 1.0425 0.7125 1.1775 0.7875 ;
        VIA 1.2300 0.5550 VIA12_square ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.0800 0.1125 1.1850 0.3375 ;
        RECT 0.6150 0.1125 1.0800 0.1875 ;
        VIA 1.1325 0.2625 VIA12_square ;
        END
    END B1
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.1125 0.4125 0.5775 0.4875 ;
        VIA 0.2400 0.4500 VIA12_square ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.1125 0.2625 0.5775 0.3375 ;
        VIA 0.4200 0.3000 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.9225 0.8625 1.3875 0.9375 ;
        RECT 0.9225 0.4125 0.9525 0.5775 ;
        RECT 0.8475 0.4125 0.9225 0.9375 ;
        VIA 0.9000 0.4950 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.6275 -0.0750 1.6800 0.0750 ;
        RECT 1.5225 -0.0750 1.6275 0.2475 ;
        RECT 0.1425 -0.0750 1.5225 0.0750 ;
        RECT 0.0675 -0.0750 0.1425 0.2550 ;
        RECT 0.0000 -0.0750 0.0675 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.6125 0.9750 1.6800 1.1250 ;
        RECT 1.5375 0.8025 1.6125 1.1250 ;
        RECT 1.2150 0.9750 1.5375 1.1250 ;
        RECT 1.0950 0.8625 1.2150 1.1250 ;
        RECT 0.0000 0.9750 1.0950 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.5450 0.1575 1.6050 0.2175 ;
        RECT 1.5450 0.8325 1.6050 0.8925 ;
        RECT 1.4475 0.4800 1.5075 0.5400 ;
        RECT 1.3350 0.8100 1.3950 0.8700 ;
        RECT 1.2300 0.4950 1.2900 0.5550 ;
        RECT 1.1250 0.8625 1.1850 0.9225 ;
        RECT 1.0275 0.4725 1.0875 0.5325 ;
        RECT 0.9150 0.1575 0.9750 0.2175 ;
        RECT 0.9150 0.8325 0.9750 0.8925 ;
        RECT 0.7050 0.1575 0.7650 0.2175 ;
        RECT 0.7050 0.8325 0.7650 0.8925 ;
        RECT 0.6000 0.4800 0.6600 0.5400 ;
        RECT 0.4950 0.6825 0.5550 0.7425 ;
        RECT 0.3900 0.4950 0.4500 0.5550 ;
        RECT 0.2850 0.8325 0.3450 0.8925 ;
        RECT 0.1800 0.4950 0.2400 0.5550 ;
        RECT 0.0750 0.1575 0.1350 0.2175 ;
        RECT 0.0750 0.7800 0.1350 0.8400 ;
        LAYER M1 ;
        RECT 1.3125 0.7125 1.4175 0.9000 ;
        RECT 1.2525 0.2850 1.3275 0.6375 ;
        RECT 1.0200 0.7125 1.3125 0.7875 ;
        RECT 1.1925 0.4725 1.2525 0.6375 ;
        RECT 1.1175 0.1800 1.1775 0.3975 ;
        RECT 1.0800 0.1800 1.1175 0.5625 ;
        RECT 1.0275 0.3300 1.0800 0.5625 ;
        RECT 0.9450 0.7125 1.0200 0.9000 ;
        RECT 0.8625 0.1500 1.0050 0.2550 ;
        RECT 0.8475 0.4125 0.9525 0.5775 ;
        RECT 0.2550 0.8250 0.9450 0.9000 ;
        RECT 0.6975 0.1500 0.8625 0.3375 ;
        RECT 0.5775 0.4575 0.8475 0.5775 ;
        RECT 0.1425 0.6750 0.8175 0.7500 ;
        RECT 0.6225 0.1500 0.6975 0.2250 ;
        RECT 0.3675 0.2175 0.4725 0.5775 ;
        RECT 0.2175 0.2100 0.2925 0.6000 ;
        RECT 0.1800 0.3675 0.2175 0.6000 ;
        RECT 0.0675 0.6750 0.1425 0.8700 ;
    END
END AOI33_1000


MACRO AOI33_1010
    CLASS CORE ;
    FOREIGN AOI33_1010 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.6800 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 0.7725 0.2625 0.8625 0.3375 ;
        RECT 0.6975 0.2625 0.7725 0.9375 ;
        RECT 0.2325 0.8625 0.6975 0.9375 ;
        VIA 0.7800 0.3000 VIA12_square ;
        VIA 0.7350 0.7125 VIA12_square ;
        END
    END ZN
    PIN B3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.5225 0.3675 1.6275 0.6825 ;
        RECT 1.4475 0.4500 1.5225 0.5700 ;
        END
    END B3
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.2750 0.7125 1.6200 0.7875 ;
        RECT 1.1700 0.4725 1.2750 0.7875 ;
        RECT 1.0425 0.7125 1.1700 0.7875 ;
        VIA 1.2225 0.5550 VIA12_square ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.0350 0.1125 1.1400 0.3375 ;
        RECT 0.6075 0.1125 1.0350 0.1875 ;
        VIA 1.0875 0.2625 VIA12_square ;
        END
    END B1
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.1125 0.4125 0.5775 0.4875 ;
        VIA 0.2400 0.4500 VIA12_square ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.1125 0.2625 0.5775 0.3375 ;
        VIA 0.4200 0.3000 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.9225 0.8625 1.3875 0.9375 ;
        RECT 0.9225 0.4125 0.9525 0.5775 ;
        RECT 0.8475 0.4125 0.9225 0.9375 ;
        VIA 0.9000 0.4950 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.6275 -0.0750 1.6800 0.0750 ;
        RECT 1.5225 -0.0750 1.6275 0.2775 ;
        RECT 0.1425 -0.0750 1.5225 0.0750 ;
        RECT 0.0675 -0.0750 0.1425 0.2550 ;
        RECT 0.0000 -0.0750 0.0675 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.6125 0.9750 1.6800 1.1250 ;
        RECT 1.5375 0.8025 1.6125 1.1250 ;
        RECT 1.2150 0.9750 1.5375 1.1250 ;
        RECT 1.0950 0.8625 1.2150 1.1250 ;
        RECT 0.0000 0.9750 1.0950 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.5450 0.1875 1.6050 0.2475 ;
        RECT 1.5450 0.8325 1.6050 0.8925 ;
        RECT 1.4475 0.4800 1.5075 0.5400 ;
        RECT 1.3350 0.7425 1.3950 0.8025 ;
        RECT 1.2300 0.4950 1.2900 0.5550 ;
        RECT 1.1250 0.8625 1.1850 0.9225 ;
        RECT 1.0275 0.4725 1.0875 0.5325 ;
        RECT 0.9150 0.1800 0.9750 0.2400 ;
        RECT 0.9150 0.8325 0.9750 0.8925 ;
        RECT 0.7050 0.2025 0.7650 0.2625 ;
        RECT 0.7050 0.8325 0.7650 0.8925 ;
        RECT 0.6000 0.4800 0.6600 0.5400 ;
        RECT 0.4950 0.6825 0.5550 0.7425 ;
        RECT 0.3900 0.4950 0.4500 0.5550 ;
        RECT 0.2850 0.8325 0.3450 0.8925 ;
        RECT 0.1800 0.4950 0.2400 0.5550 ;
        RECT 0.0750 0.1575 0.1350 0.2175 ;
        RECT 0.0750 0.7575 0.1350 0.8175 ;
        LAYER M1 ;
        RECT 1.3200 0.7125 1.4100 0.8325 ;
        RECT 1.2225 0.2850 1.3275 0.6375 ;
        RECT 1.0200 0.7125 1.3200 0.7875 ;
        RECT 1.1850 0.4725 1.2225 0.6375 ;
        RECT 1.1100 0.1800 1.1400 0.4050 ;
        RECT 1.0500 0.1800 1.1100 0.5625 ;
        RECT 1.0275 0.3300 1.0500 0.5625 ;
        RECT 0.9450 0.7125 1.0200 0.9000 ;
        RECT 0.8625 0.1500 0.9750 0.2700 ;
        RECT 0.8475 0.4125 0.9525 0.5775 ;
        RECT 0.2550 0.8250 0.9450 0.9000 ;
        RECT 0.6600 0.1500 0.8625 0.3375 ;
        RECT 0.5775 0.4575 0.8475 0.5775 ;
        RECT 0.1425 0.6750 0.8175 0.7500 ;
        RECT 0.3675 0.2175 0.4725 0.5775 ;
        RECT 0.2175 0.2100 0.2925 0.6000 ;
        RECT 0.1800 0.3675 0.2175 0.6000 ;
        RECT 0.0675 0.6750 0.1425 0.8475 ;
    END
END AOI33_1010


MACRO BUFF_0001
    CLASS CORE ;
    FOREIGN BUFF_0001 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.0500 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.9375 0.2175 1.0125 0.8325 ;
        RECT 0.9075 0.2175 0.9375 0.3825 ;
        RECT 0.9075 0.6675 0.9375 0.8325 ;
        RECT 0.5625 0.3075 0.9075 0.3825 ;
        RECT 0.5625 0.6675 0.9075 0.7425 ;
        RECT 0.4875 0.2250 0.5625 0.3825 ;
        RECT 0.4875 0.6675 0.5625 0.8175 ;
        END
    END Z
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.0525 0.4125 0.2625 0.6375 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.7950 -0.0750 1.0500 0.0750 ;
        RECT 0.6750 -0.0750 0.7950 0.2325 ;
        RECT 0.3750 -0.0750 0.6750 0.0750 ;
        RECT 0.2550 -0.0750 0.3750 0.1875 ;
        RECT 0.0000 -0.0750 0.2550 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.7875 0.9750 1.0500 1.1250 ;
        RECT 0.6825 0.8175 0.7875 1.1250 ;
        RECT 0.3750 0.9750 0.6825 1.1250 ;
        RECT 0.2550 0.8625 0.3750 1.1250 ;
        RECT 0.0000 0.9750 0.2550 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 0.9150 0.2700 0.9750 0.3300 ;
        RECT 0.9150 0.7200 0.9750 0.7800 ;
        RECT 0.8025 0.4875 0.8625 0.5475 ;
        RECT 0.7050 0.1500 0.7650 0.2100 ;
        RECT 0.7050 0.8400 0.7650 0.9000 ;
        RECT 0.6000 0.4800 0.6600 0.5400 ;
        RECT 0.4950 0.2775 0.5550 0.3375 ;
        RECT 0.4950 0.7125 0.5550 0.7725 ;
        RECT 0.3900 0.4800 0.4500 0.5400 ;
        RECT 0.2850 0.1200 0.3450 0.1800 ;
        RECT 0.2850 0.8625 0.3450 0.9225 ;
        RECT 0.1800 0.4800 0.2400 0.5400 ;
        RECT 0.0750 0.2100 0.1350 0.2700 ;
        RECT 0.0750 0.7425 0.1350 0.8025 ;
        LAYER M1 ;
        RECT 0.7575 0.4575 0.8625 0.5925 ;
        RECT 0.4125 0.4575 0.7575 0.5475 ;
        RECT 0.3375 0.2625 0.4125 0.7875 ;
        RECT 0.1575 0.2625 0.3375 0.3375 ;
        RECT 0.1575 0.7125 0.3375 0.7875 ;
        RECT 0.0525 0.1875 0.1575 0.3375 ;
        RECT 0.0525 0.7125 0.1575 0.8475 ;
    END
END BUFF_0001


MACRO BUFF_0011
    CLASS CORE ;
    FOREIGN BUFF_0011 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.8400 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.7275 0.3075 0.8025 0.7275 ;
        RECT 0.5625 0.3075 0.7275 0.3825 ;
        RECT 0.5625 0.6525 0.7275 0.7275 ;
        RECT 0.4875 0.2175 0.5625 0.3825 ;
        RECT 0.4875 0.6525 0.5625 0.8325 ;
        END
    END Z
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.0525 0.4125 0.2625 0.6375 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.7950 -0.0750 0.8400 0.0750 ;
        RECT 0.6750 -0.0750 0.7950 0.2325 ;
        RECT 0.3750 -0.0750 0.6750 0.0750 ;
        RECT 0.2550 -0.0750 0.3750 0.1800 ;
        RECT 0.0000 -0.0750 0.2550 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.7875 0.9750 0.8400 1.1250 ;
        RECT 0.6825 0.8025 0.7875 1.1250 ;
        RECT 0.3750 0.9750 0.6825 1.1250 ;
        RECT 0.2550 0.8625 0.3750 1.1250 ;
        RECT 0.0000 0.9750 0.2550 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 0.7050 0.1575 0.7650 0.2175 ;
        RECT 0.7050 0.8250 0.7650 0.8850 ;
        RECT 0.5925 0.4875 0.6525 0.5475 ;
        RECT 0.4950 0.2700 0.5550 0.3300 ;
        RECT 0.4950 0.6900 0.5550 0.7500 ;
        RECT 0.3900 0.4875 0.4500 0.5475 ;
        RECT 0.2850 0.1200 0.3450 0.1800 ;
        RECT 0.2850 0.8625 0.3450 0.9225 ;
        RECT 0.1800 0.4650 0.2400 0.5250 ;
        RECT 0.0750 0.2175 0.1350 0.2775 ;
        RECT 0.0750 0.7650 0.1350 0.8250 ;
        LAYER M1 ;
        RECT 0.4125 0.4575 0.6525 0.5775 ;
        RECT 0.3375 0.2625 0.4125 0.7875 ;
        RECT 0.1575 0.2625 0.3375 0.3375 ;
        RECT 0.1575 0.7125 0.3375 0.7875 ;
        RECT 0.0525 0.1950 0.1575 0.3375 ;
        RECT 0.0525 0.7125 0.1575 0.8475 ;
    END
END BUFF_0011


MACRO BUFF_0100
    CLASS CORE ;
    FOREIGN BUFF_0100 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.5200 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 1.7325 0.2625 1.8900 0.3825 ;
        RECT 1.7325 0.6600 1.8900 0.7800 ;
        RECT 1.4175 0.2625 1.7325 0.7800 ;
        RECT 1.2600 0.2625 1.4175 0.3825 ;
        RECT 1.2600 0.6600 1.4175 0.7800 ;
        VIA 1.7325 0.3225 VIA12_slot ;
        VIA 1.7325 0.7200 VIA12_slot ;
        VIA 1.4175 0.3225 VIA12_slot ;
        VIA 1.4175 0.7200 VIA12_slot ;
        END
    END Z
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.3525 0.4125 0.8175 0.4875 ;
        VIA 0.5250 0.4500 VIA12_square ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 2.4525 -0.0750 2.5200 0.0750 ;
        RECT 2.3775 -0.0750 2.4525 0.2925 ;
        RECT 2.0550 -0.0750 2.3775 0.0750 ;
        RECT 1.9350 -0.0750 2.0550 0.1875 ;
        RECT 1.6350 -0.0750 1.9350 0.0750 ;
        RECT 1.5150 -0.0750 1.6350 0.1875 ;
        RECT 1.2150 -0.0750 1.5150 0.0750 ;
        RECT 1.0950 -0.0750 1.2150 0.1875 ;
        RECT 0.7950 -0.0750 1.0950 0.0750 ;
        RECT 0.6750 -0.0750 0.7950 0.1875 ;
        RECT 0.3750 -0.0750 0.6750 0.0750 ;
        RECT 0.2550 -0.0750 0.3750 0.1875 ;
        RECT 0.0000 -0.0750 0.2550 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 2.4525 0.9750 2.5200 1.1250 ;
        RECT 2.3775 0.6375 2.4525 1.1250 ;
        RECT 2.0550 0.9750 2.3775 1.1250 ;
        RECT 1.9350 0.8550 2.0550 1.1250 ;
        RECT 1.6350 0.9750 1.9350 1.1250 ;
        RECT 1.5150 0.8550 1.6350 1.1250 ;
        RECT 1.2150 0.9750 1.5150 1.1250 ;
        RECT 1.0950 0.8550 1.2150 1.1250 ;
        RECT 0.7950 0.9750 1.0950 1.1250 ;
        RECT 0.6750 0.8175 0.7950 1.1250 ;
        RECT 0.3675 0.9750 0.6750 1.1250 ;
        RECT 0.2625 0.8100 0.3675 1.1250 ;
        RECT 0.0000 0.9750 0.2625 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 2.3850 0.1875 2.4450 0.2475 ;
        RECT 2.3850 0.6675 2.4450 0.7275 ;
        RECT 2.3850 0.8325 2.4450 0.8925 ;
        RECT 2.2800 0.4650 2.3400 0.5250 ;
        RECT 2.1750 0.2850 2.2350 0.3450 ;
        RECT 2.1750 0.6900 2.2350 0.7500 ;
        RECT 1.9650 0.8625 2.0250 0.9225 ;
        RECT 1.8600 0.4650 1.9200 0.5250 ;
        RECT 1.7550 0.2850 1.8150 0.3450 ;
        RECT 1.7550 0.6900 1.8150 0.7500 ;
        RECT 1.6500 0.4650 1.7100 0.5250 ;
        RECT 1.5450 0.1275 1.6050 0.1875 ;
        RECT 1.5450 0.8625 1.6050 0.9225 ;
        RECT 1.4400 0.4650 1.5000 0.5250 ;
        RECT 1.3350 0.2850 1.3950 0.3450 ;
        RECT 1.3350 0.6900 1.3950 0.7500 ;
        RECT 1.2300 0.4650 1.2900 0.5250 ;
        RECT 1.1250 0.1275 1.1850 0.1875 ;
        RECT 1.1250 0.8625 1.1850 0.9225 ;
        RECT 1.0200 0.4650 1.0800 0.5250 ;
        RECT 0.9150 0.2850 0.9750 0.3450 ;
        RECT 0.9150 0.6900 0.9750 0.7500 ;
        RECT 0.8100 0.4650 0.8700 0.5250 ;
        RECT 0.7050 0.1275 0.7650 0.1875 ;
        RECT 0.7050 0.8250 0.7650 0.8850 ;
        RECT 0.6000 0.4650 0.6600 0.5250 ;
        RECT 0.4950 0.2700 0.5550 0.3300 ;
        RECT 0.4950 0.6675 0.5550 0.7275 ;
        RECT 0.3900 0.4650 0.4500 0.5250 ;
        RECT 0.2850 0.1275 0.3450 0.1875 ;
        RECT 0.2850 0.8325 0.3450 0.8925 ;
        RECT 0.1800 0.4650 0.2400 0.5250 ;
        RECT 0.0750 0.2250 0.1350 0.2850 ;
        RECT 0.0750 0.7575 0.1350 0.8175 ;
        RECT 2.0700 0.4650 2.1300 0.5250 ;
        RECT 1.9650 0.1275 2.0250 0.1875 ;
        LAYER M1 ;
        RECT 0.8175 0.4575 2.3700 0.5325 ;
        RECT 0.8925 0.2625 2.2575 0.3825 ;
        RECT 0.8925 0.6600 2.2575 0.7800 ;
        RECT 0.7425 0.2625 0.8175 0.7350 ;
        RECT 0.1575 0.2625 0.7425 0.3375 ;
        RECT 0.1425 0.6600 0.7425 0.7350 ;
        RECT 0.5550 0.4125 0.6600 0.5625 ;
        RECT 0.1125 0.4125 0.5550 0.5325 ;
        RECT 0.0525 0.1950 0.1575 0.3375 ;
        RECT 0.0675 0.6600 0.1425 0.8700 ;
        LAYER M2 ;
        RECT 1.7625 0.2625 1.8900 0.3825 ;
        RECT 1.7625 0.6600 1.8900 0.7800 ;
        RECT 1.2600 0.2625 1.3875 0.3825 ;
        RECT 1.2600 0.6600 1.3875 0.7800 ;
    END
END BUFF_0100


MACRO BUFF_0101
    CLASS CORE ;
    FOREIGN BUFF_0101 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.5700 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 2.3625 0.2625 2.5200 0.3825 ;
        RECT 2.3625 0.6600 2.5200 0.7800 ;
        RECT 2.0475 0.2625 2.3625 0.7800 ;
        RECT 1.8900 0.2625 2.0475 0.3825 ;
        RECT 1.8900 0.6600 2.0475 0.7800 ;
        VIA 2.3625 0.3225 VIA12_slot ;
        VIA 2.3625 0.7200 VIA12_slot ;
        VIA 2.0475 0.3225 VIA12_slot ;
        VIA 2.0475 0.7200 VIA12_slot ;
        END
    END Z
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.7650 0.4125 0.8700 0.5550 ;
        RECT 0.1575 0.4125 0.7650 0.5250 ;
        RECT 0.0525 0.4125 0.1575 0.6825 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 3.5025 -0.0750 3.5700 0.0750 ;
        RECT 3.4275 -0.0750 3.5025 0.2925 ;
        RECT 3.1050 -0.0750 3.4275 0.0750 ;
        RECT 2.9850 -0.0750 3.1050 0.1875 ;
        RECT 2.6850 -0.0750 2.9850 0.0750 ;
        RECT 2.5650 -0.0750 2.6850 0.1875 ;
        RECT 2.2650 -0.0750 2.5650 0.0750 ;
        RECT 2.1450 -0.0750 2.2650 0.1875 ;
        RECT 1.8450 -0.0750 2.1450 0.0750 ;
        RECT 1.7250 -0.0750 1.8450 0.1875 ;
        RECT 1.4250 -0.0750 1.7250 0.0750 ;
        RECT 1.3050 -0.0750 1.4250 0.1875 ;
        RECT 1.0050 -0.0750 1.3050 0.0750 ;
        RECT 0.8850 -0.0750 1.0050 0.1875 ;
        RECT 0.5850 -0.0750 0.8850 0.0750 ;
        RECT 0.4650 -0.0750 0.5850 0.1875 ;
        RECT 0.1425 -0.0750 0.4650 0.0750 ;
        RECT 0.0675 -0.0750 0.1425 0.3000 ;
        RECT 0.0000 -0.0750 0.0675 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 3.5025 0.9750 3.5700 1.1250 ;
        RECT 3.4275 0.6375 3.5025 1.1250 ;
        RECT 3.1050 0.9750 3.4275 1.1250 ;
        RECT 2.9850 0.8550 3.1050 1.1250 ;
        RECT 2.6850 0.9750 2.9850 1.1250 ;
        RECT 2.5650 0.8550 2.6850 1.1250 ;
        RECT 2.2650 0.9750 2.5650 1.1250 ;
        RECT 2.1450 0.8550 2.2650 1.1250 ;
        RECT 1.8450 0.9750 2.1450 1.1250 ;
        RECT 1.7250 0.8550 1.8450 1.1250 ;
        RECT 1.4250 0.9750 1.7250 1.1250 ;
        RECT 1.3050 0.8550 1.4250 1.1250 ;
        RECT 1.0050 0.9750 1.3050 1.1250 ;
        RECT 0.8850 0.8175 1.0050 1.1250 ;
        RECT 0.5775 0.9750 0.8850 1.1250 ;
        RECT 0.4725 0.8100 0.5775 1.1250 ;
        RECT 0.1575 0.9750 0.4725 1.1250 ;
        RECT 0.0525 0.7875 0.1575 1.1250 ;
        RECT 0.0000 0.9750 0.0525 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 3.4350 0.1875 3.4950 0.2475 ;
        RECT 3.4350 0.6675 3.4950 0.7275 ;
        RECT 3.4350 0.8325 3.4950 0.8925 ;
        RECT 3.3300 0.4650 3.3900 0.5250 ;
        RECT 3.2250 0.2925 3.2850 0.3525 ;
        RECT 3.2250 0.6900 3.2850 0.7500 ;
        RECT 3.1200 0.4650 3.1800 0.5250 ;
        RECT 3.0150 0.1275 3.0750 0.1875 ;
        RECT 3.0150 0.8625 3.0750 0.9225 ;
        RECT 2.9100 0.4650 2.9700 0.5250 ;
        RECT 2.8050 0.2925 2.8650 0.3525 ;
        RECT 2.8050 0.6900 2.8650 0.7500 ;
        RECT 2.7000 0.4650 2.7600 0.5250 ;
        RECT 2.5950 0.1275 2.6550 0.1875 ;
        RECT 2.5950 0.8625 2.6550 0.9225 ;
        RECT 2.4900 0.4650 2.5500 0.5250 ;
        RECT 2.3850 0.2925 2.4450 0.3525 ;
        RECT 2.3850 0.6900 2.4450 0.7500 ;
        RECT 2.2800 0.4650 2.3400 0.5250 ;
        RECT 2.1750 0.1275 2.2350 0.1875 ;
        RECT 2.1750 0.8625 2.2350 0.9225 ;
        RECT 2.0700 0.4650 2.1300 0.5250 ;
        RECT 1.9650 0.2925 2.0250 0.3525 ;
        RECT 1.9650 0.6900 2.0250 0.7500 ;
        RECT 1.8600 0.4650 1.9200 0.5250 ;
        RECT 1.7550 0.1275 1.8150 0.1875 ;
        RECT 1.7550 0.8625 1.8150 0.9225 ;
        RECT 1.6500 0.4650 1.7100 0.5250 ;
        RECT 1.5450 0.2925 1.6050 0.3525 ;
        RECT 1.5450 0.6900 1.6050 0.7500 ;
        RECT 1.4400 0.4650 1.5000 0.5250 ;
        RECT 1.3350 0.1275 1.3950 0.1875 ;
        RECT 1.3350 0.8625 1.3950 0.9225 ;
        RECT 1.2300 0.4650 1.2900 0.5250 ;
        RECT 1.1250 0.2925 1.1850 0.3525 ;
        RECT 1.1250 0.6900 1.1850 0.7500 ;
        RECT 1.0200 0.4650 1.0800 0.5250 ;
        RECT 0.9150 0.1275 0.9750 0.1875 ;
        RECT 0.9150 0.8250 0.9750 0.8850 ;
        RECT 0.8100 0.4650 0.8700 0.5250 ;
        RECT 0.7050 0.2700 0.7650 0.3300 ;
        RECT 0.7050 0.6675 0.7650 0.7275 ;
        RECT 0.6000 0.4650 0.6600 0.5250 ;
        RECT 0.4950 0.1275 0.5550 0.1875 ;
        RECT 0.4950 0.8325 0.5550 0.8925 ;
        RECT 0.3900 0.4650 0.4500 0.5250 ;
        RECT 0.2850 0.2250 0.3450 0.2850 ;
        RECT 0.2850 0.7575 0.3450 0.8175 ;
        RECT 0.1800 0.4650 0.2400 0.5250 ;
        RECT 0.0750 0.1950 0.1350 0.2550 ;
        RECT 0.0750 0.8175 0.1350 0.8775 ;
        LAYER M1 ;
        RECT 1.0275 0.4575 3.4200 0.5325 ;
        RECT 1.1025 0.2625 3.3075 0.3825 ;
        RECT 1.1025 0.6600 3.3075 0.7800 ;
        RECT 0.9525 0.2625 1.0275 0.7350 ;
        RECT 0.3525 0.2625 0.9525 0.3375 ;
        RECT 0.3525 0.6600 0.9525 0.7350 ;
        RECT 0.2775 0.1950 0.3525 0.3375 ;
        RECT 0.2775 0.6600 0.3525 0.8700 ;
        LAYER M2 ;
        RECT 2.3925 0.2625 2.5200 0.3825 ;
        RECT 2.3925 0.6600 2.5200 0.7800 ;
        RECT 1.8900 0.2625 2.0175 0.3825 ;
        RECT 1.8900 0.6600 2.0175 0.7800 ;
    END
END BUFF_0101


MACRO BUFF_0110
    CLASS CORE ;
    FOREIGN BUFF_0110 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.8900 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 1.3125 0.2625 1.4700 0.3825 ;
        RECT 1.3125 0.6150 1.4700 0.7350 ;
        RECT 0.9975 0.2625 1.3125 0.7350 ;
        RECT 0.8400 0.2625 0.9975 0.3825 ;
        RECT 0.8400 0.6150 0.9975 0.7350 ;
        VIA 1.3125 0.3225 VIA12_slot ;
        VIA 1.3125 0.6750 VIA12_slot ;
        VIA 0.9975 0.3225 VIA12_slot ;
        VIA 0.9975 0.6750 VIA12_slot ;
        END
    END Z
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1575 0.4275 0.4500 0.5625 ;
        RECT 0.0525 0.3675 0.1575 0.6825 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.8225 -0.0750 1.8900 0.0750 ;
        RECT 1.7475 -0.0750 1.8225 0.2925 ;
        RECT 1.4250 -0.0750 1.7475 0.0750 ;
        RECT 1.3050 -0.0750 1.4250 0.1875 ;
        RECT 1.0050 -0.0750 1.3050 0.0750 ;
        RECT 0.8850 -0.0750 1.0050 0.1875 ;
        RECT 0.5850 -0.0750 0.8850 0.0750 ;
        RECT 0.4650 -0.0750 0.5850 0.1875 ;
        RECT 0.1425 -0.0750 0.4650 0.0750 ;
        RECT 0.0675 -0.0750 0.1425 0.2625 ;
        RECT 0.0000 -0.0750 0.0675 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.8225 0.9750 1.8900 1.1250 ;
        RECT 1.7475 0.6375 1.8225 1.1250 ;
        RECT 1.4175 0.9750 1.7475 1.1250 ;
        RECT 1.3125 0.8175 1.4175 1.1250 ;
        RECT 0.9975 0.9750 1.3125 1.1250 ;
        RECT 0.8925 0.8175 0.9975 1.1250 ;
        RECT 0.5850 0.9750 0.8925 1.1250 ;
        RECT 0.4650 0.8175 0.5850 1.1250 ;
        RECT 0.1425 0.9750 0.4650 1.1250 ;
        RECT 0.0675 0.7950 0.1425 1.1250 ;
        RECT 0.0000 0.9750 0.0675 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.7550 0.1875 1.8150 0.2475 ;
        RECT 1.7550 0.6675 1.8150 0.7275 ;
        RECT 1.7550 0.8325 1.8150 0.8925 ;
        RECT 1.6500 0.4650 1.7100 0.5250 ;
        RECT 1.5450 0.2850 1.6050 0.3450 ;
        RECT 1.5450 0.7575 1.6050 0.8175 ;
        RECT 1.4400 0.4650 1.5000 0.5250 ;
        RECT 1.3350 0.1275 1.3950 0.1875 ;
        RECT 1.3350 0.8475 1.3950 0.9075 ;
        RECT 1.2300 0.4650 1.2900 0.5250 ;
        RECT 1.1250 0.2850 1.1850 0.3450 ;
        RECT 1.1250 0.6450 1.1850 0.7050 ;
        RECT 1.0200 0.4650 1.0800 0.5250 ;
        RECT 0.9150 0.1275 0.9750 0.1875 ;
        RECT 0.9150 0.8475 0.9750 0.9075 ;
        RECT 0.8100 0.4650 0.8700 0.5250 ;
        RECT 0.7050 0.2850 0.7650 0.3450 ;
        RECT 0.7050 0.7575 0.7650 0.8175 ;
        RECT 0.6000 0.4650 0.6600 0.5250 ;
        RECT 0.4950 0.1275 0.5550 0.1875 ;
        RECT 0.4950 0.8250 0.5550 0.8850 ;
        RECT 0.3900 0.4650 0.4500 0.5250 ;
        RECT 0.2850 0.2250 0.3450 0.2850 ;
        RECT 0.2850 0.7575 0.3450 0.8175 ;
        RECT 0.1800 0.4650 0.2400 0.5250 ;
        RECT 0.0750 0.1725 0.1350 0.2325 ;
        RECT 0.0750 0.8250 0.1350 0.8850 ;
        LAYER M1 ;
        RECT 0.6075 0.4425 1.7400 0.5475 ;
        RECT 0.6825 0.2625 1.6275 0.3675 ;
        RECT 1.5375 0.6225 1.6125 0.8700 ;
        RECT 0.7725 0.6225 1.5375 0.7350 ;
        RECT 0.6975 0.6225 0.7725 0.8700 ;
        RECT 0.5325 0.2625 0.6075 0.7125 ;
        RECT 0.3675 0.2625 0.5325 0.3375 ;
        RECT 0.3525 0.6375 0.5325 0.7125 ;
        RECT 0.2775 0.6375 0.3525 0.8700 ;
        RECT 0.2625 0.1950 0.3675 0.3375 ;
        LAYER M2 ;
        RECT 1.3425 0.2625 1.4700 0.3825 ;
        RECT 1.3425 0.6150 1.4700 0.7350 ;
        RECT 0.8400 0.2625 0.9675 0.3825 ;
        RECT 0.8400 0.6150 0.9675 0.7350 ;
    END
END BUFF_0110


MACRO BUFF_0111
    CLASS CORE ;
    FOREIGN BUFF_0111 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.4700 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 0.7875 0.2625 1.1025 0.7500 ;
        VIA 0.9450 0.3450 VIA12_slot ;
        VIA 0.9450 0.6675 VIA12_slot ;
        END
    END Z
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1575 0.4275 0.4500 0.5625 ;
        RECT 0.0525 0.3675 0.1575 0.6825 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.4025 -0.0750 1.4700 0.0750 ;
        RECT 1.3275 -0.0750 1.4025 0.3150 ;
        RECT 1.0050 -0.0750 1.3275 0.0750 ;
        RECT 0.8850 -0.0750 1.0050 0.1950 ;
        RECT 0.5850 -0.0750 0.8850 0.0750 ;
        RECT 0.4650 -0.0750 0.5850 0.1875 ;
        RECT 0.1425 -0.0750 0.4650 0.0750 ;
        RECT 0.0675 -0.0750 0.1425 0.2625 ;
        RECT 0.0000 -0.0750 0.0675 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.4025 0.9750 1.4700 1.1250 ;
        RECT 1.3275 0.6375 1.4025 1.1250 ;
        RECT 0.9825 0.9750 1.3275 1.1250 ;
        RECT 0.9075 0.8175 0.9825 1.1250 ;
        RECT 0.5850 0.9750 0.9075 1.1250 ;
        RECT 0.4650 0.8175 0.5850 1.1250 ;
        RECT 0.1425 0.9750 0.4650 1.1250 ;
        RECT 0.0675 0.7950 0.1425 1.1250 ;
        RECT 0.0000 0.9750 0.0675 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.3350 0.2250 1.3950 0.2850 ;
        RECT 1.3350 0.6675 1.3950 0.7275 ;
        RECT 1.3350 0.8325 1.3950 0.8925 ;
        RECT 1.2300 0.4650 1.2900 0.5250 ;
        RECT 1.1250 0.2250 1.1850 0.2850 ;
        RECT 1.1250 0.7200 1.1850 0.7800 ;
        RECT 1.0200 0.4650 1.0800 0.5250 ;
        RECT 0.9150 0.1275 0.9750 0.1875 ;
        RECT 0.9150 0.8475 0.9750 0.9075 ;
        RECT 0.8100 0.4650 0.8700 0.5250 ;
        RECT 0.7050 0.2250 0.7650 0.2850 ;
        RECT 0.7050 0.7200 0.7650 0.7800 ;
        RECT 0.6000 0.4650 0.6600 0.5250 ;
        RECT 0.4950 0.1275 0.5550 0.1875 ;
        RECT 0.4950 0.8250 0.5550 0.8850 ;
        RECT 0.3900 0.4650 0.4500 0.5250 ;
        RECT 0.2850 0.2250 0.3450 0.2850 ;
        RECT 0.2850 0.7575 0.3450 0.8175 ;
        RECT 0.1800 0.4650 0.2400 0.5250 ;
        RECT 0.0750 0.1575 0.1350 0.2175 ;
        RECT 0.0750 0.8250 0.1350 0.8850 ;
        LAYER M1 ;
        RECT 0.6075 0.4575 1.3200 0.5325 ;
        RECT 0.7875 0.2925 1.1025 0.3825 ;
        RECT 0.6825 0.1950 0.7875 0.3825 ;
        RECT 0.6975 0.6225 0.7725 0.8325 ;
        RECT 0.5325 0.2625 0.6075 0.7125 ;
        RECT 0.3675 0.2625 0.5325 0.3375 ;
        RECT 0.3525 0.6375 0.5325 0.7125 ;
        RECT 0.2625 0.1950 0.3675 0.3375 ;
        RECT 0.2775 0.6375 0.3525 0.8700 ;
        RECT 1.1025 0.1950 1.2075 0.3825 ;
        RECT 1.1175 0.6225 1.1925 0.8325 ;
        RECT 0.7725 0.6225 1.1175 0.7125 ;
    END
END BUFF_0111


MACRO BUFF_1010
    CLASS CORE ;
    FOREIGN BUFF_1010 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.6300 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.5175 0.2175 0.5925 0.8325 ;
        RECT 0.4875 0.2175 0.5175 0.3825 ;
        RECT 0.4875 0.6675 0.5175 0.8325 ;
        END
    END Z
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.0525 0.4050 0.2625 0.6375 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.3750 -0.0750 0.6300 0.0750 ;
        RECT 0.2550 -0.0750 0.3750 0.1800 ;
        RECT 0.0000 -0.0750 0.2550 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.3750 0.9750 0.6300 1.1250 ;
        RECT 0.2550 0.8625 0.3750 1.1250 ;
        RECT 0.0000 0.9750 0.2550 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 0.4950 0.2775 0.5550 0.3375 ;
        RECT 0.4950 0.7275 0.5550 0.7875 ;
        RECT 0.3825 0.4950 0.4425 0.5550 ;
        RECT 0.2850 0.1200 0.3450 0.1800 ;
        RECT 0.2850 0.8625 0.3450 0.9225 ;
        RECT 0.1800 0.4650 0.2400 0.5250 ;
        RECT 0.0750 0.1725 0.1350 0.2325 ;
        RECT 0.0750 0.8175 0.1350 0.8775 ;
        LAYER M1 ;
        RECT 0.4125 0.4650 0.4425 0.5850 ;
        RECT 0.3375 0.2550 0.4125 0.7875 ;
        RECT 0.1575 0.2550 0.3375 0.3300 ;
        RECT 0.1575 0.7125 0.3375 0.7875 ;
        RECT 0.0525 0.1500 0.1575 0.3300 ;
        RECT 0.0525 0.7125 0.1575 0.9000 ;
    END
END BUFF_1010


MACRO BUFF_1100
    CLASS CORE ;
    FOREIGN BUFF_1100 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.6200 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 2.9925 0.2625 3.1500 0.3825 ;
        RECT 2.9925 0.6600 3.1500 0.7800 ;
        RECT 2.6775 0.2625 2.9925 0.7800 ;
        RECT 2.5200 0.2625 2.6775 0.3825 ;
        RECT 2.5200 0.6600 2.6775 0.7800 ;
        VIA 2.9925 0.3225 VIA12_slot ;
        VIA 2.9925 0.7200 VIA12_slot ;
        VIA 2.6775 0.3225 VIA12_slot ;
        VIA 2.6775 0.7200 VIA12_slot ;
        END
    END Z
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.4800 0.4125 0.9450 0.4875 ;
        VIA 0.7350 0.4500 VIA12_square ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 4.5525 -0.0750 4.6200 0.0750 ;
        RECT 4.4775 -0.0750 4.5525 0.2925 ;
        RECT 4.1550 -0.0750 4.4775 0.0750 ;
        RECT 4.0350 -0.0750 4.1550 0.1875 ;
        RECT 3.7350 -0.0750 4.0350 0.0750 ;
        RECT 3.6150 -0.0750 3.7350 0.1875 ;
        RECT 3.3150 -0.0750 3.6150 0.0750 ;
        RECT 3.1950 -0.0750 3.3150 0.1875 ;
        RECT 2.8950 -0.0750 3.1950 0.0750 ;
        RECT 2.7750 -0.0750 2.8950 0.1875 ;
        RECT 2.4750 -0.0750 2.7750 0.0750 ;
        RECT 2.3550 -0.0750 2.4750 0.1875 ;
        RECT 2.0550 -0.0750 2.3550 0.0750 ;
        RECT 1.9350 -0.0750 2.0550 0.1875 ;
        RECT 1.6350 -0.0750 1.9350 0.0750 ;
        RECT 1.5150 -0.0750 1.6350 0.1875 ;
        RECT 1.2150 -0.0750 1.5150 0.0750 ;
        RECT 1.0950 -0.0750 1.2150 0.1875 ;
        RECT 0.7950 -0.0750 1.0950 0.0750 ;
        RECT 0.6750 -0.0750 0.7950 0.1875 ;
        RECT 0.3750 -0.0750 0.6750 0.0750 ;
        RECT 0.2550 -0.0750 0.3750 0.1875 ;
        RECT 0.0000 -0.0750 0.2550 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 4.5525 0.9750 4.6200 1.1250 ;
        RECT 4.4775 0.6375 4.5525 1.1250 ;
        RECT 4.1550 0.9750 4.4775 1.1250 ;
        RECT 4.0350 0.8550 4.1550 1.1250 ;
        RECT 3.7350 0.9750 4.0350 1.1250 ;
        RECT 3.6150 0.8550 3.7350 1.1250 ;
        RECT 3.3150 0.9750 3.6150 1.1250 ;
        RECT 3.1950 0.8550 3.3150 1.1250 ;
        RECT 2.8950 0.9750 3.1950 1.1250 ;
        RECT 2.7750 0.8550 2.8950 1.1250 ;
        RECT 2.4750 0.9750 2.7750 1.1250 ;
        RECT 2.3550 0.8550 2.4750 1.1250 ;
        RECT 2.0550 0.9750 2.3550 1.1250 ;
        RECT 1.9350 0.8550 2.0550 1.1250 ;
        RECT 1.6350 0.9750 1.9350 1.1250 ;
        RECT 1.5150 0.8550 1.6350 1.1250 ;
        RECT 1.2150 0.9750 1.5150 1.1250 ;
        RECT 1.0950 0.8175 1.2150 1.1250 ;
        RECT 0.7950 0.9750 1.0950 1.1250 ;
        RECT 0.6750 0.8175 0.7950 1.1250 ;
        RECT 0.3675 0.9750 0.6750 1.1250 ;
        RECT 0.2625 0.8175 0.3675 1.1250 ;
        RECT 0.0000 0.9750 0.2625 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 4.4850 0.1875 4.5450 0.2475 ;
        RECT 4.4850 0.6675 4.5450 0.7275 ;
        RECT 4.4850 0.8325 4.5450 0.8925 ;
        RECT 4.3800 0.4650 4.4400 0.5250 ;
        RECT 4.2750 0.2925 4.3350 0.3525 ;
        RECT 4.2750 0.6900 4.3350 0.7500 ;
        RECT 4.1700 0.4650 4.2300 0.5250 ;
        RECT 4.0650 0.1275 4.1250 0.1875 ;
        RECT 4.0650 0.8625 4.1250 0.9225 ;
        RECT 3.9600 0.4650 4.0200 0.5250 ;
        RECT 3.8550 0.2925 3.9150 0.3525 ;
        RECT 3.8550 0.6900 3.9150 0.7500 ;
        RECT 3.7500 0.4650 3.8100 0.5250 ;
        RECT 3.6450 0.1275 3.7050 0.1875 ;
        RECT 3.6450 0.8625 3.7050 0.9225 ;
        RECT 3.5400 0.4650 3.6000 0.5250 ;
        RECT 3.4350 0.2925 3.4950 0.3525 ;
        RECT 3.4350 0.6900 3.4950 0.7500 ;
        RECT 3.3300 0.4650 3.3900 0.5250 ;
        RECT 3.2250 0.1275 3.2850 0.1875 ;
        RECT 3.2250 0.8625 3.2850 0.9225 ;
        RECT 3.1200 0.4650 3.1800 0.5250 ;
        RECT 3.0150 0.2925 3.0750 0.3525 ;
        RECT 3.0150 0.6900 3.0750 0.7500 ;
        RECT 2.9100 0.4650 2.9700 0.5250 ;
        RECT 2.8050 0.1275 2.8650 0.1875 ;
        RECT 2.8050 0.8625 2.8650 0.9225 ;
        RECT 2.7000 0.4650 2.7600 0.5250 ;
        RECT 2.5950 0.2925 2.6550 0.3525 ;
        RECT 2.5950 0.6900 2.6550 0.7500 ;
        RECT 2.4900 0.4650 2.5500 0.5250 ;
        RECT 2.3850 0.1275 2.4450 0.1875 ;
        RECT 2.3850 0.8625 2.4450 0.9225 ;
        RECT 2.2800 0.4650 2.3400 0.5250 ;
        RECT 2.1750 0.2925 2.2350 0.3525 ;
        RECT 2.1750 0.6900 2.2350 0.7500 ;
        RECT 2.0700 0.4650 2.1300 0.5250 ;
        RECT 1.9650 0.1275 2.0250 0.1875 ;
        RECT 1.9650 0.8625 2.0250 0.9225 ;
        RECT 1.8600 0.4650 1.9200 0.5250 ;
        RECT 1.7550 0.2925 1.8150 0.3525 ;
        RECT 1.7550 0.6900 1.8150 0.7500 ;
        RECT 1.6500 0.4650 1.7100 0.5250 ;
        RECT 1.5450 0.1275 1.6050 0.1875 ;
        RECT 1.5450 0.8625 1.6050 0.9225 ;
        RECT 1.4400 0.4650 1.5000 0.5250 ;
        RECT 1.3350 0.2925 1.3950 0.3525 ;
        RECT 1.3350 0.6900 1.3950 0.7500 ;
        RECT 1.2300 0.4650 1.2900 0.5250 ;
        RECT 1.1250 0.1275 1.1850 0.1875 ;
        RECT 1.1250 0.8250 1.1850 0.8850 ;
        RECT 1.0200 0.4650 1.0800 0.5250 ;
        RECT 0.9150 0.2700 0.9750 0.3300 ;
        RECT 0.9150 0.6750 0.9750 0.7350 ;
        RECT 0.8100 0.4650 0.8700 0.5250 ;
        RECT 0.7050 0.1275 0.7650 0.1875 ;
        RECT 0.7050 0.8250 0.7650 0.8850 ;
        RECT 0.6000 0.4650 0.6600 0.5250 ;
        RECT 0.4950 0.2700 0.5550 0.3300 ;
        RECT 0.4950 0.6750 0.5550 0.7350 ;
        RECT 0.3900 0.4650 0.4500 0.5250 ;
        RECT 0.2850 0.1275 0.3450 0.1875 ;
        RECT 0.2850 0.8475 0.3450 0.9075 ;
        RECT 0.1800 0.4650 0.2400 0.5250 ;
        RECT 0.0750 0.2250 0.1350 0.2850 ;
        RECT 0.0750 0.7575 0.1350 0.8175 ;
        LAYER M1 ;
        RECT 1.2375 0.4575 4.4700 0.5325 ;
        RECT 1.3125 0.2625 4.3575 0.3825 ;
        RECT 1.3125 0.6600 4.3575 0.7800 ;
        RECT 1.1625 0.2625 1.2375 0.7425 ;
        RECT 0.1425 0.2625 1.1625 0.3375 ;
        RECT 0.1425 0.6675 1.1625 0.7425 ;
        RECT 0.9750 0.4125 1.0800 0.5550 ;
        RECT 0.1125 0.4125 0.9750 0.5250 ;
        RECT 0.0675 0.1950 0.1425 0.3375 ;
        RECT 0.0675 0.6675 0.1425 0.8700 ;
        LAYER M2 ;
        RECT 3.0225 0.2625 3.1500 0.3825 ;
        RECT 3.0225 0.6600 3.1500 0.7800 ;
        RECT 2.5200 0.2625 2.6475 0.3825 ;
        RECT 2.5200 0.6600 2.6475 0.7800 ;
    END
END BUFF_1100


MACRO CKAN2_0011
    CLASS CORE ;
    FOREIGN CKAN2_0011 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.0500 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.9375 0.3075 1.0125 0.7425 ;
        RECT 0.7725 0.3075 0.9375 0.3825 ;
        RECT 0.7725 0.6675 0.9375 0.7425 ;
        RECT 0.6975 0.2175 0.7725 0.3825 ;
        RECT 0.6975 0.6675 0.7725 0.8325 ;
        END
    END Z
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.1875 0.2625 0.6525 0.3375 ;
        VIA 0.4800 0.3000 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.4275 0.8625 0.7800 0.9375 ;
        RECT 0.3525 0.4125 0.4275 0.9375 ;
        RECT 0.1875 0.4125 0.3525 0.4875 ;
        RECT 0.0675 0.8625 0.3525 0.9375 ;
        VIA 0.2700 0.4500 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.0050 -0.0750 1.0500 0.0750 ;
        RECT 0.8850 -0.0750 1.0050 0.2175 ;
        RECT 0.5925 -0.0750 0.8850 0.0750 ;
        RECT 0.4575 -0.0750 0.5925 0.1800 ;
        RECT 0.0000 -0.0750 0.4575 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.0050 0.9750 1.0500 1.1250 ;
        RECT 0.8850 0.8325 1.0050 1.1250 ;
        RECT 0.6000 0.9750 0.8850 1.1250 ;
        RECT 0.4650 0.8550 0.6000 1.1250 ;
        RECT 0.1650 0.9750 0.4650 1.1250 ;
        RECT 0.0450 0.8250 0.1650 1.1250 ;
        RECT 0.0000 0.9750 0.0450 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 0.9150 0.1575 0.9750 0.2175 ;
        RECT 0.9150 0.8325 0.9750 0.8925 ;
        RECT 0.8025 0.4950 0.8625 0.5550 ;
        RECT 0.7050 0.2625 0.7650 0.3225 ;
        RECT 0.7050 0.7275 0.7650 0.7875 ;
        RECT 0.5925 0.4950 0.6525 0.5550 ;
        RECT 0.4950 0.1200 0.5550 0.1800 ;
        RECT 0.4950 0.8550 0.5550 0.9150 ;
        RECT 0.3975 0.4800 0.4575 0.5400 ;
        RECT 0.2850 0.8175 0.3450 0.8775 ;
        RECT 0.1875 0.4800 0.2475 0.5400 ;
        RECT 0.0750 0.1575 0.1350 0.2175 ;
        RECT 0.0750 0.8325 0.1350 0.8925 ;
        LAYER M1 ;
        RECT 0.6225 0.4650 0.8625 0.5850 ;
        RECT 0.5475 0.4650 0.6225 0.7500 ;
        RECT 0.4725 0.2550 0.5625 0.3450 ;
        RECT 0.3675 0.6750 0.5475 0.7500 ;
        RECT 0.3975 0.2550 0.4725 0.5700 ;
        RECT 0.2625 0.6750 0.3675 0.9000 ;
        RECT 0.1875 0.3375 0.3225 0.6000 ;
        RECT 0.1125 0.6750 0.2625 0.7500 ;
        RECT 0.1125 0.1500 0.1650 0.2250 ;
        RECT 0.0375 0.1500 0.1125 0.7500 ;
    END
END CKAN2_0011


MACRO CKAN2_0100
    CLASS CORE ;
    FOREIGN CKAN2_0100 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.1500 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 2.3625 0.2775 2.5200 0.3975 ;
        RECT 2.3625 0.6225 2.5200 0.7425 ;
        RECT 2.0475 0.2775 2.3625 0.7425 ;
        RECT 1.8900 0.2775 2.0475 0.3975 ;
        RECT 1.8900 0.6225 2.0475 0.7425 ;
        VIA 2.3625 0.3375 VIA12_slot ;
        VIA 2.3625 0.6825 VIA12_slot ;
        VIA 2.0475 0.3375 VIA12_slot ;
        VIA 2.0475 0.6825 VIA12_slot ;
        END
    END Z
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.1850 0.4350 1.3050 0.5400 ;
        RECT 1.1100 0.4350 1.1850 0.7875 ;
        RECT 0.5625 0.7125 1.1100 0.7875 ;
        RECT 0.4875 0.4500 0.5625 0.7875 ;
        VIA 1.2225 0.4875 VIA12_square ;
        VIA 0.5250 0.5325 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.8400 0.4725 1.1100 0.5775 ;
        RECT 0.7650 0.3300 0.8400 0.5775 ;
        RECT 0.2475 0.3300 0.7650 0.4050 ;
        RECT 0.1575 0.3300 0.2475 0.5550 ;
        RECT 0.0525 0.3300 0.1575 0.6825 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 3.0975 -0.0750 3.1500 0.0750 ;
        RECT 2.9925 -0.0750 3.0975 0.3075 ;
        RECT 2.6850 -0.0750 2.9925 0.0750 ;
        RECT 2.5650 -0.0750 2.6850 0.2025 ;
        RECT 2.2650 -0.0750 2.5650 0.0750 ;
        RECT 2.1450 -0.0750 2.2650 0.2025 ;
        RECT 1.8450 -0.0750 2.1450 0.0750 ;
        RECT 1.7250 -0.0750 1.8450 0.2025 ;
        RECT 1.4100 -0.0750 1.7250 0.0750 ;
        RECT 1.3350 -0.0750 1.4100 0.2625 ;
        RECT 0.5775 -0.0750 1.3350 0.0750 ;
        RECT 0.4725 -0.0750 0.5775 0.2550 ;
        RECT 0.0000 -0.0750 0.4725 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 3.0975 0.9750 3.1500 1.1250 ;
        RECT 2.9925 0.6450 3.0975 1.1250 ;
        RECT 2.6850 0.9750 2.9925 1.1250 ;
        RECT 2.5650 0.8250 2.6850 1.1250 ;
        RECT 2.2650 0.9750 2.5650 1.1250 ;
        RECT 2.1450 0.8250 2.2650 1.1250 ;
        RECT 1.8450 0.9750 2.1450 1.1250 ;
        RECT 1.7250 0.8250 1.8450 1.1250 ;
        RECT 1.4175 0.9750 1.7250 1.1250 ;
        RECT 1.3125 0.8100 1.4175 1.1250 ;
        RECT 0.9975 0.9750 1.3125 1.1250 ;
        RECT 0.8925 0.8100 0.9975 1.1250 ;
        RECT 0.5775 0.9750 0.8925 1.1250 ;
        RECT 0.4725 0.8100 0.5775 1.1250 ;
        RECT 0.1425 0.9750 0.4725 1.1250 ;
        RECT 0.0675 0.8025 0.1425 1.1250 ;
        RECT 0.0000 0.9750 0.0675 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 3.0150 0.2175 3.0750 0.2775 ;
        RECT 3.0150 0.6675 3.0750 0.7275 ;
        RECT 3.0150 0.8325 3.0750 0.8925 ;
        RECT 2.9100 0.4800 2.9700 0.5400 ;
        RECT 2.8050 0.3075 2.8650 0.3675 ;
        RECT 2.8050 0.6525 2.8650 0.7125 ;
        RECT 2.7000 0.4800 2.7600 0.5400 ;
        RECT 2.5950 0.1350 2.6550 0.1950 ;
        RECT 2.5950 0.8325 2.6550 0.8925 ;
        RECT 2.4900 0.4800 2.5500 0.5400 ;
        RECT 2.3850 0.3075 2.4450 0.3675 ;
        RECT 2.3850 0.6525 2.4450 0.7125 ;
        RECT 2.2800 0.4800 2.3400 0.5400 ;
        RECT 2.1750 0.1350 2.2350 0.1950 ;
        RECT 2.1750 0.8325 2.2350 0.8925 ;
        RECT 2.0700 0.4800 2.1300 0.5400 ;
        RECT 1.9650 0.3075 2.0250 0.3675 ;
        RECT 1.9650 0.6525 2.0250 0.7125 ;
        RECT 1.8600 0.4800 1.9200 0.5400 ;
        RECT 1.7550 0.1350 1.8150 0.1950 ;
        RECT 1.7550 0.8325 1.8150 0.8925 ;
        RECT 1.6500 0.4800 1.7100 0.5400 ;
        RECT 1.5450 0.3075 1.6050 0.3675 ;
        RECT 1.5450 0.6525 1.6050 0.7125 ;
        RECT 1.4400 0.4800 1.5000 0.5400 ;
        RECT 1.3350 0.1725 1.3950 0.2325 ;
        RECT 1.3350 0.8325 1.3950 0.8925 ;
        RECT 1.2300 0.4800 1.2900 0.5400 ;
        RECT 1.1250 0.7950 1.1850 0.8550 ;
        RECT 1.0200 0.4950 1.0800 0.5550 ;
        RECT 0.9150 0.2325 0.9750 0.2925 ;
        RECT 0.9150 0.8325 0.9750 0.8925 ;
        RECT 0.8100 0.4950 0.8700 0.5550 ;
        RECT 0.7050 0.7950 0.7650 0.8550 ;
        RECT 0.1800 0.4650 0.2400 0.5250 ;
        RECT 0.0750 0.1725 0.1350 0.2325 ;
        RECT 0.0750 0.8325 0.1350 0.8925 ;
        RECT 0.6000 0.5025 0.6600 0.5625 ;
        RECT 0.4950 0.1725 0.5550 0.2325 ;
        RECT 0.4950 0.8325 0.5550 0.8925 ;
        RECT 0.3900 0.5025 0.4500 0.5625 ;
        RECT 0.2850 0.7950 0.3450 0.8550 ;
        LAYER M1 ;
        RECT 1.4475 0.4725 3.0000 0.5475 ;
        RECT 1.5225 0.6225 2.8950 0.7425 ;
        RECT 1.5225 0.2775 2.8875 0.3975 ;
        RECT 1.3725 0.4725 1.4475 0.7350 ;
        RECT 1.2075 0.6600 1.3725 0.7350 ;
        RECT 1.2600 0.4500 1.2975 0.5700 ;
        RECT 1.1850 0.2250 1.2600 0.5700 ;
        RECT 1.1025 0.6600 1.2075 0.8775 ;
        RECT 1.1175 0.2250 1.1850 0.3900 ;
        RECT 0.7875 0.6600 1.1025 0.7350 ;
        RECT 0.9150 0.1500 1.0425 0.3975 ;
        RECT 0.6825 0.6600 0.7875 0.8775 ;
        RECT 0.3600 0.4800 0.6900 0.5850 ;
        RECT 0.3675 0.6600 0.6825 0.7350 ;
        RECT 0.0525 0.1500 0.3975 0.2550 ;
        RECT 0.2625 0.6600 0.3675 0.8775 ;
        LAYER VIA1 ;
        RECT 1.5150 0.4725 1.5900 0.5475 ;
        RECT 0.9225 0.1950 0.9975 0.2700 ;
        RECT 0.2775 0.1650 0.3525 0.2400 ;
        LAYER M2 ;
        RECT 2.3925 0.2775 2.5200 0.3975 ;
        RECT 2.3925 0.6225 2.5200 0.7425 ;
        RECT 1.8900 0.2775 2.0175 0.3975 ;
        RECT 1.8900 0.6225 2.0175 0.7425 ;
        RECT 1.5150 0.1950 1.5900 0.5925 ;
        RECT 0.3975 0.1950 1.5150 0.2700 ;
        RECT 0.2325 0.1500 0.3975 0.2700 ;
    END
END CKAN2_0100


MACRO CKAN2_0111
    CLASS CORE ;
    FOREIGN CKAN2_0111 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.8900 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 1.2075 0.2475 1.5225 0.7650 ;
        VIA 1.3650 0.3300 VIA12_slot ;
        VIA 1.3650 0.6825 VIA12_slot ;
        END
    END Z
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.7725 0.3300 0.8775 0.5700 ;
        RECT 0.2475 0.3300 0.7725 0.4050 ;
        RECT 0.1575 0.3300 0.2475 0.5550 ;
        RECT 0.0525 0.3300 0.1575 0.6825 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.5625 0.8625 1.0275 0.9375 ;
        RECT 0.4875 0.4500 0.5625 0.9375 ;
        VIA 0.5250 0.5325 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.8375 -0.0750 1.8900 0.0750 ;
        RECT 1.7325 -0.0750 1.8375 0.3075 ;
        RECT 1.4250 -0.0750 1.7325 0.0750 ;
        RECT 1.3050 -0.0750 1.4250 0.1950 ;
        RECT 0.9975 -0.0750 1.3050 0.0750 ;
        RECT 0.8925 -0.0750 0.9975 0.2475 ;
        RECT 0.1575 -0.0750 0.8925 0.0750 ;
        RECT 0.0525 -0.0750 0.1575 0.2475 ;
        RECT 0.0000 -0.0750 0.0525 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.8375 0.9750 1.8900 1.1250 ;
        RECT 1.7325 0.6450 1.8375 1.1250 ;
        RECT 1.4250 0.9750 1.7325 1.1250 ;
        RECT 1.3050 0.8250 1.4250 1.1250 ;
        RECT 0.9975 0.9750 1.3050 1.1250 ;
        RECT 0.8925 0.8100 0.9975 1.1250 ;
        RECT 0.5775 0.9750 0.8925 1.1250 ;
        RECT 0.4725 0.8100 0.5775 1.1250 ;
        RECT 0.1425 0.9750 0.4725 1.1250 ;
        RECT 0.0675 0.8025 0.1425 1.1250 ;
        RECT 0.0000 0.9750 0.0675 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.7550 0.2175 1.8150 0.2775 ;
        RECT 1.7550 0.6675 1.8150 0.7275 ;
        RECT 1.7550 0.8325 1.8150 0.8925 ;
        RECT 1.6500 0.4725 1.7100 0.5325 ;
        RECT 1.5450 0.3000 1.6050 0.3600 ;
        RECT 1.5450 0.6525 1.6050 0.7125 ;
        RECT 1.4400 0.4725 1.5000 0.5325 ;
        RECT 1.3350 0.1275 1.3950 0.1875 ;
        RECT 1.3350 0.8325 1.3950 0.8925 ;
        RECT 1.2300 0.4725 1.2900 0.5325 ;
        RECT 1.1250 0.3000 1.1850 0.3600 ;
        RECT 1.1250 0.6525 1.1850 0.7125 ;
        RECT 1.0200 0.4725 1.0800 0.5325 ;
        RECT 0.9150 0.1650 0.9750 0.2250 ;
        RECT 0.9150 0.8325 0.9750 0.8925 ;
        RECT 0.8100 0.4800 0.8700 0.5400 ;
        RECT 0.7050 0.7800 0.7650 0.8400 ;
        RECT 0.6000 0.5025 0.6600 0.5625 ;
        RECT 0.4950 0.1725 0.5550 0.2325 ;
        RECT 0.4950 0.8325 0.5550 0.8925 ;
        RECT 0.3900 0.5025 0.4500 0.5625 ;
        RECT 0.2850 0.7800 0.3450 0.8400 ;
        RECT 0.1800 0.4650 0.2400 0.5250 ;
        RECT 0.0750 0.1650 0.1350 0.2250 ;
        RECT 0.0750 0.8325 0.1350 0.8925 ;
        LAYER M1 ;
        RECT 1.0275 0.4650 1.7700 0.5400 ;
        RECT 1.1025 0.6225 1.6350 0.7425 ;
        RECT 1.1025 0.2700 1.6275 0.3900 ;
        RECT 0.9525 0.4650 1.0275 0.7350 ;
        RECT 0.7875 0.6600 0.9525 0.7350 ;
        RECT 0.4650 0.1500 0.8175 0.2550 ;
        RECT 0.6825 0.6600 0.7875 0.8625 ;
        RECT 0.3600 0.4800 0.6900 0.5850 ;
        RECT 0.3675 0.6600 0.6825 0.7350 ;
        RECT 0.2625 0.6600 0.3675 0.8625 ;
        LAYER VIA1 ;
        RECT 0.8025 0.6600 0.8775 0.7350 ;
        RECT 0.6975 0.1800 0.7725 0.2550 ;
        LAYER M2 ;
        RECT 0.8025 0.6600 0.9225 0.7350 ;
        RECT 0.7275 0.1500 0.8025 0.7350 ;
        RECT 0.6675 0.1500 0.7275 0.2850 ;
    END
END CKAN2_0111


MACRO CKAN2_1000
    CLASS CORE ;
    FOREIGN CKAN2_1000 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.8400 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.7275 0.1500 0.8025 0.8325 ;
        RECT 0.6750 0.1500 0.7275 0.2625 ;
        RECT 0.6975 0.6675 0.7275 0.8325 ;
        END
    END Z
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.1425 0.2625 0.6075 0.3375 ;
        VIA 0.4650 0.3000 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.4800 0.8625 0.6525 0.9375 ;
        RECT 0.4050 0.4125 0.4800 0.9375 ;
        RECT 0.1725 0.4125 0.4050 0.4875 ;
        RECT 0.1125 0.8625 0.4050 0.9375 ;
        VIA 0.2550 0.4500 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.5925 -0.0750 0.8400 0.0750 ;
        RECT 0.4575 -0.0750 0.5925 0.1800 ;
        RECT 0.0000 -0.0750 0.4575 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.6000 0.9750 0.8400 1.1250 ;
        RECT 0.4500 0.8400 0.6000 1.1250 ;
        RECT 0.1650 0.9750 0.4500 1.1250 ;
        RECT 0.0450 0.8250 0.1650 1.1250 ;
        RECT 0.0000 0.9750 0.0450 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 0.7050 0.1575 0.7650 0.2175 ;
        RECT 0.7050 0.7275 0.7650 0.7875 ;
        RECT 0.5925 0.4950 0.6525 0.5550 ;
        RECT 0.4950 0.1200 0.5550 0.1800 ;
        RECT 0.4950 0.8550 0.5550 0.9150 ;
        RECT 0.3900 0.4800 0.4500 0.5400 ;
        RECT 0.2850 0.8175 0.3450 0.8775 ;
        RECT 0.1875 0.4800 0.2475 0.5400 ;
        RECT 0.0750 0.1575 0.1350 0.2175 ;
        RECT 0.0750 0.8325 0.1350 0.8925 ;
        LAYER M1 ;
        RECT 0.6225 0.4650 0.6525 0.5850 ;
        RECT 0.5475 0.4650 0.6225 0.7500 ;
        RECT 0.4575 0.2550 0.5625 0.3450 ;
        RECT 0.3675 0.6750 0.5475 0.7500 ;
        RECT 0.3825 0.2550 0.4575 0.5700 ;
        RECT 0.2625 0.6750 0.3675 0.9000 ;
        RECT 0.1875 0.3000 0.2925 0.6000 ;
        RECT 0.1125 0.6750 0.2625 0.7500 ;
        RECT 0.1125 0.1500 0.1650 0.2250 ;
        RECT 0.0375 0.1500 0.1125 0.7500 ;
    END
END CKAN2_1000


MACRO CKAN2_1010
    CLASS CORE ;
    FOREIGN CKAN2_1010 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.8400 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.7275 0.2175 0.8025 0.8325 ;
        RECT 0.6975 0.2175 0.7275 0.3825 ;
        RECT 0.6975 0.6675 0.7275 0.8325 ;
        END
    END Z
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.4575 0.2625 0.5475 0.3375 ;
        RECT 0.3750 0.2625 0.4575 0.5700 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.2250 0.1800 0.3000 0.5700 ;
        RECT 0.1875 0.4500 0.2250 0.5700 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.5925 -0.0750 0.8400 0.0750 ;
        RECT 0.4575 -0.0750 0.5925 0.1875 ;
        RECT 0.0000 -0.0750 0.4575 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.5850 0.9750 0.8400 1.1250 ;
        RECT 0.4650 0.8250 0.5850 1.1250 ;
        RECT 0.1650 0.9750 0.4650 1.1250 ;
        RECT 0.0450 0.8250 0.1650 1.1250 ;
        RECT 0.0000 0.9750 0.0450 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 0.7050 0.2625 0.7650 0.3225 ;
        RECT 0.7050 0.7275 0.7650 0.7875 ;
        RECT 0.5925 0.4950 0.6525 0.5550 ;
        RECT 0.4950 0.1275 0.5550 0.1875 ;
        RECT 0.4950 0.8250 0.5550 0.8850 ;
        RECT 0.3900 0.4800 0.4500 0.5400 ;
        RECT 0.2850 0.7875 0.3450 0.8475 ;
        RECT 0.1875 0.4800 0.2475 0.5400 ;
        RECT 0.0750 0.2400 0.1350 0.3000 ;
        RECT 0.0750 0.8325 0.1350 0.8925 ;
        LAYER M1 ;
        RECT 0.6225 0.4650 0.6525 0.5850 ;
        RECT 0.5475 0.4650 0.6225 0.7500 ;
        RECT 0.3675 0.6750 0.5475 0.7500 ;
        RECT 0.2625 0.6750 0.3675 0.8700 ;
        RECT 0.1125 0.6750 0.2625 0.7500 ;
        RECT 0.1125 0.2100 0.1425 0.3300 ;
        RECT 0.0375 0.2100 0.1125 0.7500 ;
    END
END CKAN2_1010


MACRO CKB_0000
    CLASS CORE ;
    FOREIGN CKB_0000 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.6700 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 3.6225 0.2625 3.7800 0.3825 ;
        RECT 3.6225 0.6600 3.7800 0.7800 ;
        RECT 3.3075 0.2625 3.6225 0.7800 ;
        RECT 3.1500 0.2625 3.3075 0.3825 ;
        RECT 3.1500 0.6600 3.3075 0.7800 ;
        VIA 3.6225 0.3225 VIA12_slot ;
        VIA 3.6225 0.7200 VIA12_slot ;
        VIA 3.3075 0.3225 VIA12_slot ;
        VIA 3.3075 0.7200 VIA12_slot ;
        END
    END Z
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1425 0.4275 1.2900 0.5625 ;
        RECT 0.0675 0.3675 0.1425 0.6825 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 5.6025 -0.0750 5.6700 0.0750 ;
        RECT 5.5275 -0.0750 5.6025 0.2925 ;
        RECT 5.2050 -0.0750 5.5275 0.0750 ;
        RECT 5.0850 -0.0750 5.2050 0.1875 ;
        RECT 4.7850 -0.0750 5.0850 0.0750 ;
        RECT 4.6650 -0.0750 4.7850 0.1875 ;
        RECT 4.3650 -0.0750 4.6650 0.0750 ;
        RECT 4.2450 -0.0750 4.3650 0.1875 ;
        RECT 3.9450 -0.0750 4.2450 0.0750 ;
        RECT 3.8250 -0.0750 3.9450 0.1875 ;
        RECT 3.5250 -0.0750 3.8250 0.0750 ;
        RECT 3.4050 -0.0750 3.5250 0.1875 ;
        RECT 3.1050 -0.0750 3.4050 0.0750 ;
        RECT 2.9850 -0.0750 3.1050 0.1875 ;
        RECT 2.6850 -0.0750 2.9850 0.0750 ;
        RECT 2.5650 -0.0750 2.6850 0.1875 ;
        RECT 2.2650 -0.0750 2.5650 0.0750 ;
        RECT 2.1450 -0.0750 2.2650 0.1875 ;
        RECT 1.8450 -0.0750 2.1450 0.0750 ;
        RECT 1.7250 -0.0750 1.8450 0.1875 ;
        RECT 1.4250 -0.0750 1.7250 0.0750 ;
        RECT 1.3050 -0.0750 1.4250 0.1875 ;
        RECT 1.0050 -0.0750 1.3050 0.0750 ;
        RECT 0.8850 -0.0750 1.0050 0.1875 ;
        RECT 0.5850 -0.0750 0.8850 0.0750 ;
        RECT 0.4650 -0.0750 0.5850 0.1875 ;
        RECT 0.1650 -0.0750 0.4650 0.0750 ;
        RECT 0.0450 -0.0750 0.1650 0.2700 ;
        RECT 0.0000 -0.0750 0.0450 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 5.6025 0.9750 5.6700 1.1250 ;
        RECT 5.5275 0.6375 5.6025 1.1250 ;
        RECT 5.2050 0.9750 5.5275 1.1250 ;
        RECT 5.0850 0.8550 5.2050 1.1250 ;
        RECT 4.7850 0.9750 5.0850 1.1250 ;
        RECT 4.6650 0.8550 4.7850 1.1250 ;
        RECT 4.3650 0.9750 4.6650 1.1250 ;
        RECT 4.2450 0.8550 4.3650 1.1250 ;
        RECT 3.9450 0.9750 4.2450 1.1250 ;
        RECT 3.8250 0.8550 3.9450 1.1250 ;
        RECT 3.5250 0.9750 3.8250 1.1250 ;
        RECT 3.4050 0.8550 3.5250 1.1250 ;
        RECT 3.1050 0.9750 3.4050 1.1250 ;
        RECT 2.9850 0.8550 3.1050 1.1250 ;
        RECT 2.6850 0.9750 2.9850 1.1250 ;
        RECT 2.5650 0.8550 2.6850 1.1250 ;
        RECT 2.2650 0.9750 2.5650 1.1250 ;
        RECT 2.1450 0.8550 2.2650 1.1250 ;
        RECT 1.8450 0.9750 2.1450 1.1250 ;
        RECT 1.7250 0.8550 1.8450 1.1250 ;
        RECT 1.4250 0.9750 1.7250 1.1250 ;
        RECT 1.3050 0.8175 1.4250 1.1250 ;
        RECT 1.0050 0.9750 1.3050 1.1250 ;
        RECT 0.8850 0.8175 1.0050 1.1250 ;
        RECT 0.5850 0.9750 0.8850 1.1250 ;
        RECT 0.4650 0.8175 0.5850 1.1250 ;
        RECT 0.1575 0.9750 0.4650 1.1250 ;
        RECT 0.0525 0.8100 0.1575 1.1250 ;
        RECT 0.0000 0.9750 0.0525 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 5.5350 0.1875 5.5950 0.2475 ;
        RECT 5.5350 0.6675 5.5950 0.7275 ;
        RECT 5.5350 0.8325 5.5950 0.8925 ;
        RECT 5.4300 0.4650 5.4900 0.5250 ;
        RECT 5.3250 0.2925 5.3850 0.3525 ;
        RECT 5.3250 0.6900 5.3850 0.7500 ;
        RECT 5.2200 0.4650 5.2800 0.5250 ;
        RECT 5.1150 0.1275 5.1750 0.1875 ;
        RECT 5.1150 0.8625 5.1750 0.9225 ;
        RECT 5.0100 0.4650 5.0700 0.5250 ;
        RECT 4.9050 0.2925 4.9650 0.3525 ;
        RECT 4.9050 0.6900 4.9650 0.7500 ;
        RECT 4.8000 0.4650 4.8600 0.5250 ;
        RECT 4.6950 0.1275 4.7550 0.1875 ;
        RECT 4.6950 0.8625 4.7550 0.9225 ;
        RECT 4.5900 0.4650 4.6500 0.5250 ;
        RECT 4.4850 0.2925 4.5450 0.3525 ;
        RECT 4.4850 0.6900 4.5450 0.7500 ;
        RECT 4.3800 0.4650 4.4400 0.5250 ;
        RECT 4.2750 0.1275 4.3350 0.1875 ;
        RECT 4.2750 0.8625 4.3350 0.9225 ;
        RECT 4.1700 0.4650 4.2300 0.5250 ;
        RECT 4.0650 0.2925 4.1250 0.3525 ;
        RECT 4.0650 0.6900 4.1250 0.7500 ;
        RECT 3.9600 0.4650 4.0200 0.5250 ;
        RECT 3.8550 0.1275 3.9150 0.1875 ;
        RECT 3.8550 0.8625 3.9150 0.9225 ;
        RECT 3.7500 0.4650 3.8100 0.5250 ;
        RECT 3.6450 0.2925 3.7050 0.3525 ;
        RECT 3.6450 0.6900 3.7050 0.7500 ;
        RECT 3.5400 0.4650 3.6000 0.5250 ;
        RECT 3.4350 0.1275 3.4950 0.1875 ;
        RECT 3.4350 0.8625 3.4950 0.9225 ;
        RECT 3.3300 0.4650 3.3900 0.5250 ;
        RECT 3.2250 0.2925 3.2850 0.3525 ;
        RECT 3.2250 0.6900 3.2850 0.7500 ;
        RECT 3.1200 0.4650 3.1800 0.5250 ;
        RECT 3.0150 0.1275 3.0750 0.1875 ;
        RECT 3.0150 0.8625 3.0750 0.9225 ;
        RECT 2.9100 0.4650 2.9700 0.5250 ;
        RECT 2.8050 0.2925 2.8650 0.3525 ;
        RECT 2.8050 0.6900 2.8650 0.7500 ;
        RECT 2.7000 0.4650 2.7600 0.5250 ;
        RECT 2.5950 0.1275 2.6550 0.1875 ;
        RECT 2.5950 0.8625 2.6550 0.9225 ;
        RECT 2.4900 0.4650 2.5500 0.5250 ;
        RECT 2.3850 0.2925 2.4450 0.3525 ;
        RECT 2.3850 0.6900 2.4450 0.7500 ;
        RECT 2.2800 0.4650 2.3400 0.5250 ;
        RECT 2.1750 0.1275 2.2350 0.1875 ;
        RECT 2.1750 0.8625 2.2350 0.9225 ;
        RECT 2.0700 0.4650 2.1300 0.5250 ;
        RECT 1.9650 0.2925 2.0250 0.3525 ;
        RECT 1.9650 0.6900 2.0250 0.7500 ;
        RECT 1.8600 0.4650 1.9200 0.5250 ;
        RECT 1.7550 0.1275 1.8150 0.1875 ;
        RECT 1.7550 0.8625 1.8150 0.9225 ;
        RECT 1.6500 0.4650 1.7100 0.5250 ;
        RECT 1.5450 0.2925 1.6050 0.3525 ;
        RECT 1.5450 0.6900 1.6050 0.7500 ;
        RECT 1.4400 0.4650 1.5000 0.5250 ;
        RECT 1.3350 0.1275 1.3950 0.1875 ;
        RECT 1.3350 0.8250 1.3950 0.8850 ;
        RECT 1.2300 0.4650 1.2900 0.5250 ;
        RECT 1.1250 0.2700 1.1850 0.3300 ;
        RECT 1.1250 0.6750 1.1850 0.7350 ;
        RECT 1.0200 0.4650 1.0800 0.5250 ;
        RECT 0.9150 0.1275 0.9750 0.1875 ;
        RECT 0.9150 0.8250 0.9750 0.8850 ;
        RECT 0.8100 0.4650 0.8700 0.5250 ;
        RECT 0.7050 0.2700 0.7650 0.3300 ;
        RECT 0.7050 0.6750 0.7650 0.7350 ;
        RECT 0.6000 0.4650 0.6600 0.5250 ;
        RECT 0.4950 0.1275 0.5550 0.1875 ;
        RECT 0.4950 0.8250 0.5550 0.8850 ;
        RECT 0.3900 0.4650 0.4500 0.5250 ;
        RECT 0.2850 0.2250 0.3450 0.2850 ;
        RECT 0.2850 0.7575 0.3450 0.8175 ;
        RECT 0.1800 0.4650 0.2400 0.5250 ;
        RECT 0.0750 0.1950 0.1350 0.2550 ;
        RECT 0.0750 0.8325 0.1350 0.8925 ;
        LAYER M1 ;
        RECT 1.4475 0.4575 5.5200 0.5325 ;
        RECT 1.5225 0.2625 5.4075 0.3825 ;
        RECT 1.5225 0.6600 5.4075 0.7800 ;
        RECT 1.3725 0.2625 1.4475 0.7425 ;
        RECT 0.3675 0.2625 1.3725 0.3375 ;
        RECT 0.3525 0.6675 1.3725 0.7425 ;
        RECT 0.2625 0.1950 0.3675 0.3375 ;
        RECT 0.2775 0.6675 0.3525 0.8700 ;
        LAYER M2 ;
        RECT 3.6525 0.2625 3.7800 0.3825 ;
        RECT 3.6525 0.6600 3.7800 0.7800 ;
        RECT 3.1500 0.2625 3.2775 0.3825 ;
        RECT 3.1500 0.6600 3.2775 0.7800 ;
    END
END CKB_0000


MACRO CKB_0001
    CLASS CORE ;
    FOREIGN CKB_0001 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.0500 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.9375 0.3000 1.0125 0.7275 ;
        RECT 0.5625 0.3000 0.9375 0.3750 ;
        RECT 0.5625 0.6525 0.9375 0.7275 ;
        RECT 0.4875 0.2175 0.5625 0.3750 ;
        RECT 0.4875 0.6525 0.5625 0.8325 ;
        END
    END Z
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.0975 0.4125 0.5625 0.4875 ;
        VIA 0.1800 0.4500 VIA12_square ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.7950 -0.0750 1.0500 0.0750 ;
        RECT 0.6750 -0.0750 0.7950 0.2250 ;
        RECT 0.3750 -0.0750 0.6750 0.0750 ;
        RECT 0.2550 -0.0750 0.3750 0.1800 ;
        RECT 0.0000 -0.0750 0.2550 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.7875 0.9750 1.0500 1.1250 ;
        RECT 0.6825 0.8025 0.7875 1.1250 ;
        RECT 0.3675 0.9750 0.6825 1.1250 ;
        RECT 0.2625 0.8400 0.3675 1.1250 ;
        RECT 0.0000 0.9750 0.2625 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 0.9150 0.3075 0.9750 0.3675 ;
        RECT 0.9150 0.6600 0.9750 0.7200 ;
        RECT 0.8025 0.4875 0.8625 0.5475 ;
        RECT 0.7050 0.1500 0.7650 0.2100 ;
        RECT 0.7050 0.8250 0.7650 0.8850 ;
        RECT 0.6000 0.4875 0.6600 0.5475 ;
        RECT 0.4950 0.2700 0.5550 0.3300 ;
        RECT 0.4950 0.6900 0.5550 0.7500 ;
        RECT 0.3900 0.4875 0.4500 0.5475 ;
        RECT 0.2850 0.1200 0.3450 0.1800 ;
        RECT 0.2850 0.8625 0.3450 0.9225 ;
        RECT 0.1800 0.4875 0.2400 0.5475 ;
        RECT 0.0750 0.2175 0.1350 0.2775 ;
        RECT 0.0750 0.7650 0.1350 0.8250 ;
        LAYER M1 ;
        RECT 0.4125 0.4575 0.8625 0.5775 ;
        RECT 0.3375 0.2625 0.4125 0.7650 ;
        RECT 0.1575 0.2625 0.3375 0.3375 ;
        RECT 0.1575 0.6900 0.3375 0.7650 ;
        RECT 0.0525 0.4125 0.2625 0.6075 ;
        RECT 0.0525 0.1950 0.1575 0.3375 ;
        RECT 0.0525 0.6900 0.1575 0.8475 ;
    END
END CKB_0001


MACRO CKB_0011
    CLASS CORE ;
    FOREIGN CKB_0011 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.8400 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.7275 0.3075 0.8025 0.7275 ;
        RECT 0.5625 0.3075 0.7275 0.3825 ;
        RECT 0.5625 0.6525 0.7275 0.7275 ;
        RECT 0.4875 0.2175 0.5625 0.3825 ;
        RECT 0.4875 0.6525 0.5625 0.8325 ;
        END
    END Z
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.0975 0.4125 0.5625 0.4875 ;
        VIA 0.1800 0.4500 VIA12_square ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.7950 -0.0750 0.8400 0.0750 ;
        RECT 0.6750 -0.0750 0.7950 0.2325 ;
        RECT 0.3750 -0.0750 0.6750 0.0750 ;
        RECT 0.2550 -0.0750 0.3750 0.1800 ;
        RECT 0.0000 -0.0750 0.2550 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.7875 0.9750 0.8400 1.1250 ;
        RECT 0.6825 0.8025 0.7875 1.1250 ;
        RECT 0.3675 0.9750 0.6825 1.1250 ;
        RECT 0.2625 0.8400 0.3675 1.1250 ;
        RECT 0.0000 0.9750 0.2625 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 0.7050 0.1575 0.7650 0.2175 ;
        RECT 0.7050 0.8250 0.7650 0.8850 ;
        RECT 0.5925 0.4875 0.6525 0.5475 ;
        RECT 0.4950 0.2700 0.5550 0.3300 ;
        RECT 0.4950 0.6900 0.5550 0.7500 ;
        RECT 0.3900 0.4875 0.4500 0.5475 ;
        RECT 0.2850 0.1200 0.3450 0.1800 ;
        RECT 0.2850 0.8625 0.3450 0.9225 ;
        RECT 0.1800 0.4650 0.2400 0.5250 ;
        RECT 0.0750 0.2175 0.1350 0.2775 ;
        RECT 0.0750 0.7650 0.1350 0.8250 ;
        LAYER M1 ;
        RECT 0.4125 0.4575 0.6525 0.5775 ;
        RECT 0.3375 0.2625 0.4125 0.7650 ;
        RECT 0.1575 0.2625 0.3375 0.3375 ;
        RECT 0.1575 0.6900 0.3375 0.7650 ;
        RECT 0.0525 0.4125 0.2625 0.6075 ;
        RECT 0.0525 0.1950 0.1575 0.3375 ;
        RECT 0.0525 0.6900 0.1575 0.8475 ;
    END
END CKB_0011


MACRO CKB_0100
    CLASS CORE ;
    FOREIGN CKB_0100 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.5200 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 1.7325 0.2625 1.8900 0.3825 ;
        RECT 1.7325 0.6600 1.8900 0.7800 ;
        RECT 1.4175 0.2625 1.7325 0.7800 ;
        RECT 1.2600 0.2625 1.4175 0.3825 ;
        RECT 1.2600 0.6600 1.4175 0.7800 ;
        VIA 1.7325 0.3225 VIA12_slot ;
        VIA 1.7325 0.7200 VIA12_slot ;
        VIA 1.4175 0.3225 VIA12_slot ;
        VIA 1.4175 0.7200 VIA12_slot ;
        END
    END Z
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.6450 0.4125 1.1100 0.4875 ;
        RECT 0.4800 0.4125 0.6450 0.5175 ;
        VIA 0.5625 0.4650 VIA12_square ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 2.4525 -0.0750 2.5200 0.0750 ;
        RECT 2.3775 -0.0750 2.4525 0.2925 ;
        RECT 2.0550 -0.0750 2.3775 0.0750 ;
        RECT 1.9350 -0.0750 2.0550 0.1875 ;
        RECT 1.6350 -0.0750 1.9350 0.0750 ;
        RECT 1.5150 -0.0750 1.6350 0.1875 ;
        RECT 1.2150 -0.0750 1.5150 0.0750 ;
        RECT 1.0950 -0.0750 1.2150 0.1875 ;
        RECT 0.7950 -0.0750 1.0950 0.0750 ;
        RECT 0.6750 -0.0750 0.7950 0.1875 ;
        RECT 0.3750 -0.0750 0.6750 0.0750 ;
        RECT 0.2550 -0.0750 0.3750 0.1875 ;
        RECT 0.0000 -0.0750 0.2550 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 2.4525 0.9750 2.5200 1.1250 ;
        RECT 2.3775 0.6375 2.4525 1.1250 ;
        RECT 2.0550 0.9750 2.3775 1.1250 ;
        RECT 1.9350 0.8550 2.0550 1.1250 ;
        RECT 1.6350 0.9750 1.9350 1.1250 ;
        RECT 1.5150 0.8550 1.6350 1.1250 ;
        RECT 1.2150 0.9750 1.5150 1.1250 ;
        RECT 1.0950 0.8550 1.2150 1.1250 ;
        RECT 0.7950 0.9750 1.0950 1.1250 ;
        RECT 0.6750 0.8175 0.7950 1.1250 ;
        RECT 0.3675 0.9750 0.6750 1.1250 ;
        RECT 0.2625 0.8100 0.3675 1.1250 ;
        RECT 0.0000 0.9750 0.2625 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 2.3850 0.1875 2.4450 0.2475 ;
        RECT 2.3850 0.6675 2.4450 0.7275 ;
        RECT 2.3850 0.8325 2.4450 0.8925 ;
        RECT 2.2800 0.4650 2.3400 0.5250 ;
        RECT 2.1750 0.2850 2.2350 0.3450 ;
        RECT 2.1750 0.6900 2.2350 0.7500 ;
        RECT 1.9650 0.1275 2.0250 0.1875 ;
        RECT 1.9650 0.8625 2.0250 0.9225 ;
        RECT 1.8600 0.4650 1.9200 0.5250 ;
        RECT 1.7550 0.2850 1.8150 0.3450 ;
        RECT 1.7550 0.6900 1.8150 0.7500 ;
        RECT 1.6500 0.4650 1.7100 0.5250 ;
        RECT 1.5450 0.1275 1.6050 0.1875 ;
        RECT 1.5450 0.8625 1.6050 0.9225 ;
        RECT 1.4400 0.4650 1.5000 0.5250 ;
        RECT 1.3350 0.2850 1.3950 0.3450 ;
        RECT 1.3350 0.6900 1.3950 0.7500 ;
        RECT 1.2300 0.4650 1.2900 0.5250 ;
        RECT 1.1250 0.1275 1.1850 0.1875 ;
        RECT 1.1250 0.8625 1.1850 0.9225 ;
        RECT 1.0200 0.4650 1.0800 0.5250 ;
        RECT 0.9150 0.2850 0.9750 0.3450 ;
        RECT 0.9150 0.6900 0.9750 0.7500 ;
        RECT 0.8100 0.4650 0.8700 0.5250 ;
        RECT 0.7050 0.1275 0.7650 0.1875 ;
        RECT 0.7050 0.8250 0.7650 0.8850 ;
        RECT 0.6000 0.4650 0.6600 0.5250 ;
        RECT 0.4950 0.2700 0.5550 0.3300 ;
        RECT 0.4950 0.6675 0.5550 0.7275 ;
        RECT 0.3900 0.4650 0.4500 0.5250 ;
        RECT 0.2850 0.1275 0.3450 0.1875 ;
        RECT 0.2850 0.8325 0.3450 0.8925 ;
        RECT 0.1800 0.4650 0.2400 0.5250 ;
        RECT 0.0750 0.2250 0.1350 0.2850 ;
        RECT 0.0750 0.7575 0.1350 0.8175 ;
        RECT 2.0700 0.4650 2.1300 0.5250 ;
        LAYER M1 ;
        RECT 0.8175 0.4575 2.3700 0.5325 ;
        RECT 0.8925 0.2625 2.2575 0.3825 ;
        RECT 0.8925 0.6600 2.2575 0.7800 ;
        RECT 0.7425 0.2625 0.8175 0.7350 ;
        RECT 0.1575 0.2625 0.7425 0.3375 ;
        RECT 0.1425 0.6600 0.7425 0.7350 ;
        RECT 0.1125 0.4275 0.6600 0.5625 ;
        RECT 0.0525 0.1950 0.1575 0.3375 ;
        RECT 0.0675 0.6600 0.1425 0.8700 ;
        LAYER M2 ;
        RECT 1.7625 0.2625 1.8900 0.3825 ;
        RECT 1.7625 0.6600 1.8900 0.7800 ;
        RECT 1.2600 0.2625 1.3875 0.3825 ;
        RECT 1.2600 0.6600 1.3875 0.7800 ;
    END
END CKB_0100


MACRO CKB_0101
    CLASS CORE ;
    FOREIGN CKB_0101 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.5700 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 2.3625 0.2625 2.5200 0.3825 ;
        RECT 2.3625 0.6600 2.5200 0.7800 ;
        RECT 2.0475 0.2625 2.3625 0.7800 ;
        RECT 1.8900 0.2625 2.0475 0.3825 ;
        RECT 1.8900 0.6600 2.0475 0.7800 ;
        VIA 2.3625 0.3225 VIA12_slot ;
        VIA 2.3625 0.7200 VIA12_slot ;
        VIA 2.0475 0.3225 VIA12_slot ;
        VIA 2.0475 0.7200 VIA12_slot ;
        END
    END Z
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1425 0.4275 0.8700 0.5625 ;
        RECT 0.0675 0.3675 0.1425 0.6825 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 3.5250 -0.0750 3.5700 0.0750 ;
        RECT 3.4050 -0.0750 3.5250 0.2925 ;
        RECT 3.1050 -0.0750 3.4050 0.0750 ;
        RECT 2.9850 -0.0750 3.1050 0.1875 ;
        RECT 2.6850 -0.0750 2.9850 0.0750 ;
        RECT 2.5650 -0.0750 2.6850 0.1875 ;
        RECT 2.2650 -0.0750 2.5650 0.0750 ;
        RECT 2.1450 -0.0750 2.2650 0.1875 ;
        RECT 1.8450 -0.0750 2.1450 0.0750 ;
        RECT 1.7250 -0.0750 1.8450 0.1875 ;
        RECT 1.4250 -0.0750 1.7250 0.0750 ;
        RECT 1.3050 -0.0750 1.4250 0.1875 ;
        RECT 1.0050 -0.0750 1.3050 0.0750 ;
        RECT 0.8850 -0.0750 1.0050 0.1875 ;
        RECT 0.5850 -0.0750 0.8850 0.0750 ;
        RECT 0.4650 -0.0750 0.5850 0.1875 ;
        RECT 0.1575 -0.0750 0.4650 0.0750 ;
        RECT 0.0525 -0.0750 0.1575 0.2475 ;
        RECT 0.0000 -0.0750 0.0525 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 3.5250 0.9750 3.5700 1.1250 ;
        RECT 3.4050 0.6375 3.5250 1.1250 ;
        RECT 3.1050 0.9750 3.4050 1.1250 ;
        RECT 2.9850 0.8550 3.1050 1.1250 ;
        RECT 2.6850 0.9750 2.9850 1.1250 ;
        RECT 2.5650 0.8550 2.6850 1.1250 ;
        RECT 2.2650 0.9750 2.5650 1.1250 ;
        RECT 2.1450 0.8550 2.2650 1.1250 ;
        RECT 1.8450 0.9750 2.1450 1.1250 ;
        RECT 1.7250 0.8550 1.8450 1.1250 ;
        RECT 1.4250 0.9750 1.7250 1.1250 ;
        RECT 1.3050 0.8550 1.4250 1.1250 ;
        RECT 1.0050 0.9750 1.3050 1.1250 ;
        RECT 0.8850 0.8175 1.0050 1.1250 ;
        RECT 0.5775 0.9750 0.8850 1.1250 ;
        RECT 0.4725 0.8100 0.5775 1.1250 ;
        RECT 0.1575 0.9750 0.4725 1.1250 ;
        RECT 0.0525 0.8025 0.1575 1.1250 ;
        RECT 0.0000 0.9750 0.0525 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 3.4350 0.1875 3.4950 0.2475 ;
        RECT 3.4350 0.6675 3.4950 0.7275 ;
        RECT 3.4350 0.8325 3.4950 0.8925 ;
        RECT 3.3300 0.4650 3.3900 0.5250 ;
        RECT 3.2250 0.2925 3.2850 0.3525 ;
        RECT 3.2250 0.6900 3.2850 0.7500 ;
        RECT 3.1200 0.4650 3.1800 0.5250 ;
        RECT 3.0150 0.1275 3.0750 0.1875 ;
        RECT 3.0150 0.8625 3.0750 0.9225 ;
        RECT 2.9100 0.4650 2.9700 0.5250 ;
        RECT 2.8050 0.2925 2.8650 0.3525 ;
        RECT 2.8050 0.6900 2.8650 0.7500 ;
        RECT 2.7000 0.4650 2.7600 0.5250 ;
        RECT 2.5950 0.1275 2.6550 0.1875 ;
        RECT 2.5950 0.8625 2.6550 0.9225 ;
        RECT 2.4900 0.4650 2.5500 0.5250 ;
        RECT 2.3850 0.2925 2.4450 0.3525 ;
        RECT 2.3850 0.6900 2.4450 0.7500 ;
        RECT 2.2800 0.4650 2.3400 0.5250 ;
        RECT 2.1750 0.1275 2.2350 0.1875 ;
        RECT 2.1750 0.8625 2.2350 0.9225 ;
        RECT 2.0700 0.4650 2.1300 0.5250 ;
        RECT 1.9650 0.2925 2.0250 0.3525 ;
        RECT 1.9650 0.6900 2.0250 0.7500 ;
        RECT 1.8600 0.4650 1.9200 0.5250 ;
        RECT 1.7550 0.1275 1.8150 0.1875 ;
        RECT 1.7550 0.8625 1.8150 0.9225 ;
        RECT 1.6500 0.4650 1.7100 0.5250 ;
        RECT 1.5450 0.2925 1.6050 0.3525 ;
        RECT 1.5450 0.6900 1.6050 0.7500 ;
        RECT 1.4400 0.4650 1.5000 0.5250 ;
        RECT 1.3350 0.1275 1.3950 0.1875 ;
        RECT 1.3350 0.8625 1.3950 0.9225 ;
        RECT 1.2300 0.4650 1.2900 0.5250 ;
        RECT 1.1250 0.2925 1.1850 0.3525 ;
        RECT 1.1250 0.6900 1.1850 0.7500 ;
        RECT 1.0200 0.4650 1.0800 0.5250 ;
        RECT 0.9150 0.1275 0.9750 0.1875 ;
        RECT 0.9150 0.8250 0.9750 0.8850 ;
        RECT 0.8100 0.4650 0.8700 0.5250 ;
        RECT 0.7050 0.2700 0.7650 0.3300 ;
        RECT 0.7050 0.6675 0.7650 0.7275 ;
        RECT 0.6000 0.4650 0.6600 0.5250 ;
        RECT 0.4950 0.1275 0.5550 0.1875 ;
        RECT 0.4950 0.8325 0.5550 0.8925 ;
        RECT 0.3900 0.4650 0.4500 0.5250 ;
        RECT 0.2850 0.2250 0.3450 0.2850 ;
        RECT 0.2850 0.7050 0.3450 0.7650 ;
        RECT 0.1800 0.4650 0.2400 0.5250 ;
        RECT 0.0750 0.1575 0.1350 0.2175 ;
        RECT 0.0750 0.8325 0.1350 0.8925 ;
        LAYER M1 ;
        RECT 1.0275 0.4575 3.4200 0.5325 ;
        RECT 1.1025 0.2625 3.3075 0.3825 ;
        RECT 1.1025 0.6600 3.3075 0.7800 ;
        RECT 0.9525 0.2625 1.0275 0.7350 ;
        RECT 0.3525 0.2625 0.9525 0.3375 ;
        RECT 0.3525 0.6600 0.9525 0.7350 ;
        RECT 0.2775 0.1950 0.3525 0.3375 ;
        RECT 0.2775 0.6600 0.3525 0.8100 ;
        LAYER M2 ;
        RECT 2.3925 0.2625 2.5200 0.3825 ;
        RECT 2.3925 0.6600 2.5200 0.7800 ;
        RECT 1.8900 0.2625 2.0175 0.3825 ;
        RECT 1.8900 0.6600 2.0175 0.7800 ;
    END
END CKB_0101


MACRO CKB_0110
    CLASS CORE ;
    FOREIGN CKB_0110 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.8900 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 1.3125 0.2850 1.4700 0.4050 ;
        RECT 1.3125 0.6075 1.4700 0.7275 ;
        RECT 0.9975 0.2850 1.3125 0.7275 ;
        RECT 0.8400 0.2850 0.9975 0.4050 ;
        RECT 0.8400 0.6075 0.9975 0.7275 ;
        VIA 1.3125 0.3450 VIA12_slot ;
        VIA 1.3125 0.6675 VIA12_slot ;
        VIA 0.9975 0.3450 VIA12_slot ;
        VIA 0.9975 0.6675 VIA12_slot ;
        END
    END Z
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1575 0.4275 0.4500 0.5625 ;
        RECT 0.0525 0.3525 0.1575 0.6825 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.8225 -0.0750 1.8900 0.0750 ;
        RECT 1.7475 -0.0750 1.8225 0.2925 ;
        RECT 1.4250 -0.0750 1.7475 0.0750 ;
        RECT 1.3050 -0.0750 1.4250 0.1950 ;
        RECT 1.0050 -0.0750 1.3050 0.0750 ;
        RECT 0.8850 -0.0750 1.0050 0.1950 ;
        RECT 0.5850 -0.0750 0.8850 0.0750 ;
        RECT 0.4650 -0.0750 0.5850 0.1875 ;
        RECT 0.1425 -0.0750 0.4650 0.0750 ;
        RECT 0.0675 -0.0750 0.1425 0.2475 ;
        RECT 0.0000 -0.0750 0.0675 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.8375 0.9750 1.8900 1.1250 ;
        RECT 1.7325 0.6450 1.8375 1.1250 ;
        RECT 1.4025 0.9750 1.7325 1.1250 ;
        RECT 1.3275 0.8175 1.4025 1.1250 ;
        RECT 0.9825 0.9750 1.3275 1.1250 ;
        RECT 0.9075 0.8175 0.9825 1.1250 ;
        RECT 0.5850 0.9750 0.9075 1.1250 ;
        RECT 0.4650 0.8175 0.5850 1.1250 ;
        RECT 0.1425 0.9750 0.4650 1.1250 ;
        RECT 0.0675 0.7950 0.1425 1.1250 ;
        RECT 0.0000 0.9750 0.0675 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.7550 0.1875 1.8150 0.2475 ;
        RECT 1.6500 0.4725 1.7100 0.5325 ;
        RECT 1.5450 0.2250 1.6050 0.2850 ;
        RECT 1.5450 0.7575 1.6050 0.8175 ;
        RECT 1.4400 0.4725 1.5000 0.5325 ;
        RECT 1.3350 0.1275 1.3950 0.1875 ;
        RECT 1.3350 0.8475 1.3950 0.9075 ;
        RECT 1.2300 0.4725 1.2900 0.5325 ;
        RECT 1.1250 0.3000 1.1850 0.3600 ;
        RECT 1.1250 0.7575 1.1850 0.8175 ;
        RECT 1.0200 0.4725 1.0800 0.5325 ;
        RECT 0.9150 0.1275 0.9750 0.1875 ;
        RECT 0.9150 0.8475 0.9750 0.9075 ;
        RECT 0.8100 0.4725 0.8700 0.5325 ;
        RECT 0.7050 0.2250 0.7650 0.2850 ;
        RECT 0.7050 0.7575 0.7650 0.8175 ;
        RECT 0.6000 0.4725 0.6600 0.5325 ;
        RECT 0.4950 0.1275 0.5550 0.1875 ;
        RECT 0.4950 0.8250 0.5550 0.8850 ;
        RECT 0.3900 0.4650 0.4500 0.5250 ;
        RECT 0.2850 0.2250 0.3450 0.2850 ;
        RECT 0.2850 0.7575 0.3450 0.8175 ;
        RECT 0.1800 0.4650 0.2400 0.5250 ;
        RECT 0.0750 0.1575 0.1350 0.2175 ;
        RECT 0.0750 0.8250 0.1350 0.8850 ;
        RECT 1.7550 0.6675 1.8150 0.7275 ;
        RECT 1.7550 0.8325 1.8150 0.8925 ;
        LAYER M1 ;
        RECT 0.6075 0.4650 1.7400 0.5400 ;
        RECT 1.5225 0.1950 1.6275 0.3900 ;
        RECT 1.5375 0.6225 1.6125 0.8700 ;
        RECT 1.1925 0.6225 1.5375 0.7125 ;
        RECT 0.7875 0.3000 1.5225 0.3900 ;
        RECT 1.1175 0.6225 1.1925 0.8700 ;
        RECT 0.7725 0.6225 1.1175 0.7125 ;
        RECT 0.6825 0.1950 0.7875 0.3900 ;
        RECT 0.6975 0.6225 0.7725 0.8700 ;
        RECT 0.5325 0.2625 0.6075 0.7125 ;
        RECT 0.3675 0.2625 0.5325 0.3375 ;
        RECT 0.3525 0.6375 0.5325 0.7125 ;
        RECT 0.2625 0.1950 0.3675 0.3375 ;
        RECT 0.2775 0.6375 0.3525 0.8700 ;
        LAYER M2 ;
        RECT 1.3425 0.2850 1.4700 0.4050 ;
        RECT 1.3425 0.6075 1.4700 0.7275 ;
        RECT 0.8400 0.2850 0.9675 0.4050 ;
        RECT 0.8400 0.6075 0.9675 0.7275 ;
    END
END CKB_0110


MACRO CKB_0111
    CLASS CORE ;
    FOREIGN CKB_0111 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.4700 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 0.7875 0.2625 1.1025 0.7500 ;
        VIA 0.9450 0.3450 VIA12_slot ;
        VIA 0.9450 0.6675 VIA12_slot ;
        END
    END Z
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1575 0.4275 0.4500 0.5625 ;
        RECT 0.0525 0.3675 0.1575 0.6825 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.4025 -0.0750 1.4700 0.0750 ;
        RECT 1.3275 -0.0750 1.4025 0.3150 ;
        RECT 1.0050 -0.0750 1.3275 0.0750 ;
        RECT 0.8850 -0.0750 1.0050 0.1950 ;
        RECT 0.5850 -0.0750 0.8850 0.0750 ;
        RECT 0.4650 -0.0750 0.5850 0.1875 ;
        RECT 0.1425 -0.0750 0.4650 0.0750 ;
        RECT 0.0675 -0.0750 0.1425 0.2625 ;
        RECT 0.0000 -0.0750 0.0675 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.4025 0.9750 1.4700 1.1250 ;
        RECT 1.3275 0.6375 1.4025 1.1250 ;
        RECT 0.9825 0.9750 1.3275 1.1250 ;
        RECT 0.9075 0.8175 0.9825 1.1250 ;
        RECT 0.5850 0.9750 0.9075 1.1250 ;
        RECT 0.4650 0.8175 0.5850 1.1250 ;
        RECT 0.1425 0.9750 0.4650 1.1250 ;
        RECT 0.0675 0.7950 0.1425 1.1250 ;
        RECT 0.0000 0.9750 0.0675 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.3350 0.2250 1.3950 0.2850 ;
        RECT 1.3350 0.6675 1.3950 0.7275 ;
        RECT 1.3350 0.8325 1.3950 0.8925 ;
        RECT 1.2300 0.4800 1.2900 0.5400 ;
        RECT 1.1250 0.2250 1.1850 0.2850 ;
        RECT 1.1250 0.7575 1.1850 0.8175 ;
        RECT 1.0200 0.4800 1.0800 0.5400 ;
        RECT 0.9150 0.1275 0.9750 0.1875 ;
        RECT 0.9150 0.8475 0.9750 0.9075 ;
        RECT 0.8100 0.4800 0.8700 0.5400 ;
        RECT 0.7050 0.2250 0.7650 0.2850 ;
        RECT 0.7050 0.7575 0.7650 0.8175 ;
        RECT 0.6000 0.4800 0.6600 0.5400 ;
        RECT 0.4950 0.1275 0.5550 0.1875 ;
        RECT 0.4950 0.8250 0.5550 0.8850 ;
        RECT 0.3900 0.4650 0.4500 0.5250 ;
        RECT 0.2850 0.2250 0.3450 0.2850 ;
        RECT 0.2850 0.7575 0.3450 0.8175 ;
        RECT 0.1800 0.4650 0.2400 0.5250 ;
        RECT 0.0750 0.1725 0.1350 0.2325 ;
        RECT 0.0750 0.8250 0.1350 0.8850 ;
        LAYER M1 ;
        RECT 0.6075 0.4725 1.3200 0.5475 ;
        RECT 0.7875 0.3000 1.1025 0.3900 ;
        RECT 0.6825 0.1950 0.7875 0.3900 ;
        RECT 0.6975 0.6225 0.7725 0.8700 ;
        RECT 0.5325 0.2625 0.6075 0.7125 ;
        RECT 0.3675 0.2625 0.5325 0.3375 ;
        RECT 0.3525 0.6375 0.5325 0.7125 ;
        RECT 0.2625 0.1950 0.3675 0.3375 ;
        RECT 0.2775 0.6375 0.3525 0.8700 ;
        RECT 1.1025 0.1950 1.2075 0.3900 ;
        RECT 1.1175 0.6225 1.1925 0.8700 ;
        RECT 0.7725 0.6225 1.1175 0.7125 ;
    END
END CKB_0111


MACRO CKB_1000
    CLASS CORE ;
    FOREIGN CKB_1000 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.6300 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.5175 0.1500 0.5925 0.9000 ;
        RECT 0.4875 0.1500 0.5175 0.2700 ;
        RECT 0.4875 0.6675 0.5175 0.9000 ;
        END
    END Z
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.0900 0.4125 0.5550 0.4875 ;
        VIA 0.1725 0.4500 VIA12_square ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.3750 -0.0750 0.6300 0.0750 ;
        RECT 0.2550 -0.0750 0.3750 0.1875 ;
        RECT 0.0000 -0.0750 0.2550 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.3750 0.9750 0.6300 1.1250 ;
        RECT 0.2550 0.7950 0.3750 1.1250 ;
        RECT 0.0000 0.9750 0.2550 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 0.4950 0.1800 0.5550 0.2400 ;
        RECT 0.4950 0.8100 0.5550 0.8700 ;
        RECT 0.3825 0.4950 0.4425 0.5550 ;
        RECT 0.2850 0.1275 0.3450 0.1875 ;
        RECT 0.2850 0.8175 0.3450 0.8775 ;
        RECT 0.1800 0.4650 0.2400 0.5250 ;
        RECT 0.0750 0.1650 0.1350 0.2250 ;
        RECT 0.0750 0.8175 0.1350 0.8775 ;
        LAYER M1 ;
        RECT 0.4125 0.4650 0.4425 0.5850 ;
        RECT 0.3375 0.2625 0.4125 0.7125 ;
        RECT 0.1650 0.2625 0.3375 0.3375 ;
        RECT 0.1575 0.6375 0.3375 0.7125 ;
        RECT 0.0525 0.4125 0.2625 0.5625 ;
        RECT 0.0450 0.1500 0.1650 0.3375 ;
        RECT 0.0525 0.6375 0.1575 0.9000 ;
    END
END CKB_1000


MACRO CKB_1010
    CLASS CORE ;
    FOREIGN CKB_1010 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.6300 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.5175 0.1800 0.5925 0.8325 ;
        RECT 0.4950 0.1800 0.5175 0.3825 ;
        RECT 0.4950 0.6675 0.5175 0.8325 ;
        END
    END Z
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.2625 0.6375 0.4125 0.7875 ;
        RECT 0.2475 0.4425 0.2625 0.7875 ;
        RECT 0.1875 0.4425 0.2475 0.7125 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.3750 -0.0750 0.6300 0.0750 ;
        RECT 0.2550 -0.0750 0.3750 0.1875 ;
        RECT 0.0000 -0.0750 0.2550 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.3750 0.9750 0.6300 1.1250 ;
        RECT 0.2550 0.8625 0.3750 1.1250 ;
        RECT 0.0000 0.9750 0.2550 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 0.4950 0.2325 0.5550 0.2925 ;
        RECT 0.4950 0.7275 0.5550 0.7875 ;
        RECT 0.3825 0.4725 0.4425 0.5325 ;
        RECT 0.2850 0.1275 0.3450 0.1875 ;
        RECT 0.2850 0.8625 0.3450 0.9225 ;
        RECT 0.1875 0.4875 0.2475 0.5475 ;
        RECT 0.0750 0.1725 0.1350 0.2325 ;
        RECT 0.0750 0.8175 0.1350 0.8775 ;
        LAYER M1 ;
        RECT 0.4200 0.4425 0.4425 0.5625 ;
        RECT 0.3375 0.2625 0.4200 0.5625 ;
        RECT 0.1575 0.2625 0.3375 0.3375 ;
        RECT 0.1125 0.1500 0.1575 0.3375 ;
        RECT 0.1125 0.7950 0.1575 0.9000 ;
        RECT 0.0375 0.1500 0.1125 0.9000 ;
    END
END CKB_1010


MACRO CKB_1100
    CLASS CORE ;
    FOREIGN CKB_1100 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.6200 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 2.9925 0.2625 3.1500 0.3825 ;
        RECT 2.9925 0.6600 3.1500 0.7800 ;
        RECT 2.6775 0.2625 2.9925 0.7800 ;
        RECT 2.5200 0.2625 2.6775 0.3825 ;
        RECT 2.5200 0.6600 2.6775 0.7800 ;
        VIA 2.9925 0.3225 VIA12_slot ;
        VIA 2.9925 0.7200 VIA12_slot ;
        VIA 2.6775 0.3225 VIA12_slot ;
        VIA 2.6775 0.7200 VIA12_slot ;
        END
    END Z
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.0425 0.4125 1.5300 0.4875 ;
        RECT 0.8775 0.4125 1.0425 0.5175 ;
        VIA 0.9600 0.4650 VIA12_square ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 4.5525 -0.0750 4.6200 0.0750 ;
        RECT 4.4775 -0.0750 4.5525 0.2925 ;
        RECT 4.1550 -0.0750 4.4775 0.0750 ;
        RECT 4.0350 -0.0750 4.1550 0.1875 ;
        RECT 3.7350 -0.0750 4.0350 0.0750 ;
        RECT 3.6150 -0.0750 3.7350 0.1875 ;
        RECT 3.3150 -0.0750 3.6150 0.0750 ;
        RECT 3.1950 -0.0750 3.3150 0.1875 ;
        RECT 2.8950 -0.0750 3.1950 0.0750 ;
        RECT 2.7750 -0.0750 2.8950 0.1875 ;
        RECT 2.4750 -0.0750 2.7750 0.0750 ;
        RECT 2.3550 -0.0750 2.4750 0.1875 ;
        RECT 2.0550 -0.0750 2.3550 0.0750 ;
        RECT 1.9350 -0.0750 2.0550 0.1875 ;
        RECT 1.6350 -0.0750 1.9350 0.0750 ;
        RECT 1.5150 -0.0750 1.6350 0.1875 ;
        RECT 1.2150 -0.0750 1.5150 0.0750 ;
        RECT 1.0950 -0.0750 1.2150 0.1875 ;
        RECT 0.7950 -0.0750 1.0950 0.0750 ;
        RECT 0.6750 -0.0750 0.7950 0.1875 ;
        RECT 0.3750 -0.0750 0.6750 0.0750 ;
        RECT 0.2550 -0.0750 0.3750 0.1875 ;
        RECT 0.0000 -0.0750 0.2550 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 4.5525 0.9750 4.6200 1.1250 ;
        RECT 4.4775 0.6375 4.5525 1.1250 ;
        RECT 4.1550 0.9750 4.4775 1.1250 ;
        RECT 4.0350 0.8550 4.1550 1.1250 ;
        RECT 3.7350 0.9750 4.0350 1.1250 ;
        RECT 3.6150 0.8550 3.7350 1.1250 ;
        RECT 3.3150 0.9750 3.6150 1.1250 ;
        RECT 3.1950 0.8550 3.3150 1.1250 ;
        RECT 2.8950 0.9750 3.1950 1.1250 ;
        RECT 2.7750 0.8550 2.8950 1.1250 ;
        RECT 2.4750 0.9750 2.7750 1.1250 ;
        RECT 2.3550 0.8550 2.4750 1.1250 ;
        RECT 2.0550 0.9750 2.3550 1.1250 ;
        RECT 1.9350 0.8550 2.0550 1.1250 ;
        RECT 1.6350 0.9750 1.9350 1.1250 ;
        RECT 1.5150 0.8550 1.6350 1.1250 ;
        RECT 1.2150 0.9750 1.5150 1.1250 ;
        RECT 1.0950 0.8175 1.2150 1.1250 ;
        RECT 0.7950 0.9750 1.0950 1.1250 ;
        RECT 0.6750 0.8175 0.7950 1.1250 ;
        RECT 0.3675 0.9750 0.6750 1.1250 ;
        RECT 0.2625 0.8175 0.3675 1.1250 ;
        RECT 0.0000 0.9750 0.2625 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 4.4850 0.1875 4.5450 0.2475 ;
        RECT 4.4850 0.6675 4.5450 0.7275 ;
        RECT 4.4850 0.8325 4.5450 0.8925 ;
        RECT 4.3800 0.4650 4.4400 0.5250 ;
        RECT 4.2750 0.2925 4.3350 0.3525 ;
        RECT 4.2750 0.6900 4.3350 0.7500 ;
        RECT 4.1700 0.4650 4.2300 0.5250 ;
        RECT 4.0650 0.1275 4.1250 0.1875 ;
        RECT 4.0650 0.8625 4.1250 0.9225 ;
        RECT 3.9600 0.4650 4.0200 0.5250 ;
        RECT 3.8550 0.2925 3.9150 0.3525 ;
        RECT 3.8550 0.6900 3.9150 0.7500 ;
        RECT 3.7500 0.4650 3.8100 0.5250 ;
        RECT 3.6450 0.1275 3.7050 0.1875 ;
        RECT 3.6450 0.8625 3.7050 0.9225 ;
        RECT 3.5400 0.4650 3.6000 0.5250 ;
        RECT 3.4350 0.2925 3.4950 0.3525 ;
        RECT 3.4350 0.6900 3.4950 0.7500 ;
        RECT 3.3300 0.4650 3.3900 0.5250 ;
        RECT 3.2250 0.1275 3.2850 0.1875 ;
        RECT 3.2250 0.8625 3.2850 0.9225 ;
        RECT 3.1200 0.4650 3.1800 0.5250 ;
        RECT 3.0150 0.2925 3.0750 0.3525 ;
        RECT 3.0150 0.6900 3.0750 0.7500 ;
        RECT 2.9100 0.4650 2.9700 0.5250 ;
        RECT 2.8050 0.1275 2.8650 0.1875 ;
        RECT 2.8050 0.8625 2.8650 0.9225 ;
        RECT 2.7000 0.4650 2.7600 0.5250 ;
        RECT 2.5950 0.2925 2.6550 0.3525 ;
        RECT 2.5950 0.6900 2.6550 0.7500 ;
        RECT 2.4900 0.4650 2.5500 0.5250 ;
        RECT 2.3850 0.1275 2.4450 0.1875 ;
        RECT 2.3850 0.8625 2.4450 0.9225 ;
        RECT 2.2800 0.4650 2.3400 0.5250 ;
        RECT 2.1750 0.2925 2.2350 0.3525 ;
        RECT 2.1750 0.6900 2.2350 0.7500 ;
        RECT 2.0700 0.4650 2.1300 0.5250 ;
        RECT 1.9650 0.1275 2.0250 0.1875 ;
        RECT 1.9650 0.8625 2.0250 0.9225 ;
        RECT 1.8600 0.4650 1.9200 0.5250 ;
        RECT 1.7550 0.2925 1.8150 0.3525 ;
        RECT 1.7550 0.6900 1.8150 0.7500 ;
        RECT 1.6500 0.4650 1.7100 0.5250 ;
        RECT 1.5450 0.1275 1.6050 0.1875 ;
        RECT 1.5450 0.8625 1.6050 0.9225 ;
        RECT 1.4400 0.4650 1.5000 0.5250 ;
        RECT 1.3350 0.2925 1.3950 0.3525 ;
        RECT 1.3350 0.6900 1.3950 0.7500 ;
        RECT 1.2300 0.4650 1.2900 0.5250 ;
        RECT 1.1250 0.1275 1.1850 0.1875 ;
        RECT 1.1250 0.8250 1.1850 0.8850 ;
        RECT 1.0200 0.4650 1.0800 0.5250 ;
        RECT 0.9150 0.2700 0.9750 0.3300 ;
        RECT 0.9150 0.6750 0.9750 0.7350 ;
        RECT 0.8100 0.4650 0.8700 0.5250 ;
        RECT 0.7050 0.1275 0.7650 0.1875 ;
        RECT 0.7050 0.8250 0.7650 0.8850 ;
        RECT 0.6000 0.4650 0.6600 0.5250 ;
        RECT 0.4950 0.2700 0.5550 0.3300 ;
        RECT 0.4950 0.6750 0.5550 0.7350 ;
        RECT 0.3900 0.4650 0.4500 0.5250 ;
        RECT 0.2850 0.1275 0.3450 0.1875 ;
        RECT 0.2850 0.8475 0.3450 0.9075 ;
        RECT 0.1800 0.4650 0.2400 0.5250 ;
        RECT 0.0750 0.2250 0.1350 0.2850 ;
        RECT 0.0750 0.7575 0.1350 0.8175 ;
        LAYER M1 ;
        RECT 1.2375 0.4575 4.4700 0.5325 ;
        RECT 1.3125 0.2625 4.3575 0.3825 ;
        RECT 1.3125 0.6600 4.3575 0.7800 ;
        RECT 1.1625 0.2625 1.2375 0.7425 ;
        RECT 0.1425 0.2625 1.1625 0.3375 ;
        RECT 0.1425 0.6675 1.1625 0.7425 ;
        RECT 0.1125 0.4275 1.0800 0.5625 ;
        RECT 0.0675 0.1950 0.1425 0.3375 ;
        RECT 0.0675 0.6675 0.1425 0.8700 ;
        LAYER M2 ;
        RECT 3.0225 0.2625 3.1500 0.3825 ;
        RECT 3.0225 0.6600 3.1500 0.7800 ;
        RECT 2.5200 0.2625 2.6475 0.3825 ;
        RECT 2.5200 0.6600 2.6475 0.7800 ;
    END
END CKB_1100


MACRO CKLNQ_0001
    CLASS CORE ;
    FOREIGN CKLNQ_0001 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.5700 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN TE
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.0900 0.7125 0.5700 0.7875 ;
        VIA 0.3150 0.7500 VIA12_square ;
        END
    END TE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 3.4575 0.3000 3.5325 0.7500 ;
        RECT 3.0825 0.3000 3.4575 0.3825 ;
        RECT 3.0825 0.6675 3.4575 0.7500 ;
        RECT 3.0075 0.2175 3.0825 0.3825 ;
        RECT 3.0075 0.6675 3.0825 0.8325 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.4275 0.2625 0.8925 0.3375 ;
        RECT 0.3525 0.2625 0.4275 0.5400 ;
        VIA 0.3900 0.4575 VIA12_square ;
        END
    END E
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 2.0250 0.4125 2.5500 0.4875 ;
        VIA 2.3100 0.4500 VIA12_square ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 3.3150 -0.0750 3.5700 0.0750 ;
        RECT 3.1950 -0.0750 3.3150 0.2250 ;
        RECT 2.8950 -0.0750 3.1950 0.0750 ;
        RECT 2.7750 -0.0750 2.8950 0.1800 ;
        RECT 2.0550 -0.0750 2.7750 0.0750 ;
        RECT 1.9350 -0.0750 2.0550 0.1875 ;
        RECT 1.4250 -0.0750 1.9350 0.0750 ;
        RECT 1.3050 -0.0750 1.4250 0.2100 ;
        RECT 0.3750 -0.0750 1.3050 0.0750 ;
        RECT 0.2550 -0.0750 0.3750 0.1800 ;
        RECT 0.0000 -0.0750 0.2550 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 3.3150 0.9750 3.5700 1.1250 ;
        RECT 3.1950 0.8250 3.3150 1.1250 ;
        RECT 2.8950 0.9750 3.1950 1.1250 ;
        RECT 2.7750 0.8700 2.8950 1.1250 ;
        RECT 2.4750 0.9750 2.7750 1.1250 ;
        RECT 2.3700 0.8025 2.4750 1.1250 ;
        RECT 2.0550 0.9750 2.3700 1.1250 ;
        RECT 1.9350 0.8625 2.0550 1.1250 ;
        RECT 1.4100 0.9750 1.9350 1.1250 ;
        RECT 1.3350 0.8400 1.4100 1.1250 ;
        RECT 0.1650 0.9750 1.3350 1.1250 ;
        RECT 0.0450 0.8250 0.1650 1.1250 ;
        RECT 0.0000 0.9750 0.0450 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 3.4350 0.3000 3.4950 0.3600 ;
        RECT 3.4350 0.6825 3.4950 0.7425 ;
        RECT 3.3225 0.4875 3.3825 0.5475 ;
        RECT 3.2250 0.1575 3.2850 0.2175 ;
        RECT 3.2250 0.8325 3.2850 0.8925 ;
        RECT 3.1200 0.4875 3.1800 0.5475 ;
        RECT 3.0150 0.2475 3.0750 0.3075 ;
        RECT 3.0150 0.7425 3.0750 0.8025 ;
        RECT 2.9100 0.4875 2.9700 0.5475 ;
        RECT 2.8050 0.1200 2.8650 0.1800 ;
        RECT 2.8050 0.8700 2.8650 0.9300 ;
        RECT 2.7000 0.4875 2.7600 0.5475 ;
        RECT 2.5950 0.8100 2.6550 0.8700 ;
        RECT 2.4900 0.4725 2.5500 0.5325 ;
        RECT 2.3850 0.2250 2.4450 0.2850 ;
        RECT 2.3850 0.8325 2.4450 0.8925 ;
        RECT 2.1750 0.2700 2.2350 0.3300 ;
        RECT 2.1750 0.7200 2.2350 0.7800 ;
        RECT 2.0700 0.4725 2.1300 0.5325 ;
        RECT 1.9650 0.1200 2.0250 0.1800 ;
        RECT 1.9650 0.8625 2.0250 0.9225 ;
        RECT 1.8675 0.4650 1.9275 0.5250 ;
        RECT 1.7550 0.2325 1.8150 0.2925 ;
        RECT 1.7550 0.6525 1.8150 0.7125 ;
        RECT 1.5450 0.1575 1.6050 0.2175 ;
        RECT 1.5450 0.8325 1.6050 0.8925 ;
        RECT 1.4325 0.6450 1.4925 0.7050 ;
        RECT 1.3350 0.1275 1.3950 0.1875 ;
        RECT 1.3350 0.8700 1.3950 0.9300 ;
        RECT 1.2300 0.3150 1.2900 0.3750 ;
        RECT 1.0200 0.3525 1.0800 0.4125 ;
        RECT 1.0200 0.6150 1.0800 0.6750 ;
        RECT 0.9150 0.1575 0.9750 0.2175 ;
        RECT 0.9150 0.8325 0.9750 0.8925 ;
        RECT 0.8175 0.3975 0.8775 0.4575 ;
        RECT 0.7050 0.1575 0.7650 0.2175 ;
        RECT 0.7050 0.8100 0.7650 0.8700 ;
        RECT 0.6075 0.5775 0.6675 0.6375 ;
        RECT 0.4950 0.2100 0.5550 0.2700 ;
        RECT 0.4950 0.8100 0.5550 0.8700 ;
        RECT 0.3900 0.4650 0.4500 0.5250 ;
        RECT 0.2850 0.1200 0.3450 0.1800 ;
        RECT 0.1725 0.4650 0.2325 0.5250 ;
        RECT 0.0750 0.2100 0.1350 0.2700 ;
        RECT 0.0750 0.8325 0.1350 0.8925 ;
        LAYER M1 ;
        RECT 2.9325 0.4575 3.3825 0.5775 ;
        RECT 2.8575 0.2550 2.9325 0.7950 ;
        RECT 2.4525 0.2550 2.8575 0.3300 ;
        RECT 2.6775 0.7200 2.8575 0.7950 ;
        RECT 2.6250 0.4050 2.7825 0.6450 ;
        RECT 2.5725 0.7200 2.6775 0.8925 ;
        RECT 2.3925 0.4425 2.5500 0.5625 ;
        RECT 2.3775 0.1800 2.4525 0.3300 ;
        RECT 2.2275 0.4125 2.3925 0.5625 ;
        RECT 1.9950 0.2625 2.2650 0.3375 ;
        RECT 1.9950 0.7125 2.2650 0.7875 ;
        RECT 2.0700 0.4425 2.2275 0.5625 ;
        RECT 1.9200 0.2625 1.9950 0.7875 ;
        RECT 1.8675 0.4350 1.9200 0.5550 ;
        RECT 1.7925 0.2025 1.8375 0.3225 ;
        RECT 1.7925 0.6300 1.8375 0.7350 ;
        RECT 1.7175 0.2025 1.7925 0.7350 ;
        RECT 1.5675 0.1500 1.6425 0.9000 ;
        RECT 1.5150 0.1500 1.5675 0.3600 ;
        RECT 1.5150 0.8250 1.5675 0.9000 ;
        RECT 1.2975 0.2850 1.5150 0.3600 ;
        RECT 1.2600 0.6150 1.4925 0.7350 ;
        RECT 1.2225 0.2850 1.2975 0.4050 ;
        RECT 1.1850 0.6150 1.2600 0.9000 ;
        RECT 0.8850 0.8100 1.1850 0.9000 ;
        RECT 1.0200 0.3225 1.1400 0.4875 ;
        RECT 0.9150 0.5625 1.0800 0.7050 ;
        RECT 0.8175 0.3675 1.0200 0.4875 ;
        RECT 0.7425 0.1500 1.0125 0.2250 ;
        RECT 0.6975 0.6150 0.9150 0.7050 ;
        RECT 0.4875 0.7800 0.7800 0.9000 ;
        RECT 0.6675 0.1500 0.7425 0.5025 ;
        RECT 0.5775 0.5775 0.6975 0.7050 ;
        RECT 0.5775 0.4125 0.6675 0.5025 ;
        RECT 0.4875 0.1800 0.5625 0.3300 ;
        RECT 0.1425 0.2550 0.4875 0.3300 ;
        RECT 0.3075 0.4050 0.4725 0.6000 ;
        RECT 0.2475 0.6750 0.3825 0.8175 ;
        RECT 0.2325 0.6750 0.2475 0.7500 ;
        RECT 0.1575 0.4350 0.2325 0.7500 ;
        RECT 0.0675 0.1800 0.1425 0.3300 ;
        LAYER VIA1 ;
        RECT 2.6775 0.5250 2.7525 0.6000 ;
        RECT 1.9200 0.5625 1.9950 0.6375 ;
        RECT 1.7175 0.3675 1.7925 0.4425 ;
        RECT 1.5675 0.7125 1.6425 0.7875 ;
        RECT 1.1850 0.7125 1.2600 0.7875 ;
        RECT 1.0650 0.3675 1.1400 0.4425 ;
        RECT 0.9600 0.5625 1.0350 0.6375 ;
        RECT 0.6225 0.4275 0.6975 0.5025 ;
        LAYER M2 ;
        RECT 2.6775 0.4800 2.7525 0.7875 ;
        RECT 1.5225 0.7125 2.6775 0.7875 ;
        RECT 0.9150 0.5625 2.0400 0.6375 ;
        RECT 1.0200 0.3675 1.8375 0.4425 ;
        RECT 0.7650 0.7125 1.3050 0.7875 ;
        RECT 0.6900 0.4275 0.7650 0.7875 ;
        RECT 0.5775 0.4275 0.6900 0.5025 ;
    END
END CKLNQ_0001


MACRO CKLNQ_0011
    CLASS CORE ;
    FOREIGN CKLNQ_0011 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.3600 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN TE
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.0900 0.7125 0.5700 0.7875 ;
        VIA 0.3150 0.7500 VIA12_square ;
        END
    END TE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 3.2475 0.3075 3.3225 0.7500 ;
        RECT 3.0825 0.3075 3.2475 0.3825 ;
        RECT 3.0825 0.6675 3.2475 0.7500 ;
        RECT 3.0075 0.2175 3.0825 0.3825 ;
        RECT 3.0075 0.6675 3.0825 0.8325 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.4275 0.2625 0.8925 0.3375 ;
        RECT 0.3525 0.2625 0.4275 0.5400 ;
        VIA 0.3900 0.4575 VIA12_square ;
        END
    END E
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 2.0250 0.4125 2.5500 0.4875 ;
        VIA 2.3100 0.4500 VIA12_square ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 3.3150 -0.0750 3.3600 0.0750 ;
        RECT 3.1950 -0.0750 3.3150 0.2250 ;
        RECT 2.8950 -0.0750 3.1950 0.0750 ;
        RECT 2.7750 -0.0750 2.8950 0.1800 ;
        RECT 2.0550 -0.0750 2.7750 0.0750 ;
        RECT 1.9350 -0.0750 2.0550 0.1875 ;
        RECT 1.4250 -0.0750 1.9350 0.0750 ;
        RECT 1.3050 -0.0750 1.4250 0.2100 ;
        RECT 0.3750 -0.0750 1.3050 0.0750 ;
        RECT 0.2550 -0.0750 0.3750 0.1800 ;
        RECT 0.0000 -0.0750 0.2550 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 3.3150 0.9750 3.3600 1.1250 ;
        RECT 3.1950 0.8250 3.3150 1.1250 ;
        RECT 2.8950 0.9750 3.1950 1.1250 ;
        RECT 2.7750 0.8700 2.8950 1.1250 ;
        RECT 2.4750 0.9750 2.7750 1.1250 ;
        RECT 2.3700 0.8025 2.4750 1.1250 ;
        RECT 2.0550 0.9750 2.3700 1.1250 ;
        RECT 1.9350 0.8625 2.0550 1.1250 ;
        RECT 1.4100 0.9750 1.9350 1.1250 ;
        RECT 1.3350 0.8400 1.4100 1.1250 ;
        RECT 0.1650 0.9750 1.3350 1.1250 ;
        RECT 0.0450 0.8250 0.1650 1.1250 ;
        RECT 0.0000 0.9750 0.0450 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 3.2250 0.1575 3.2850 0.2175 ;
        RECT 3.2250 0.8325 3.2850 0.8925 ;
        RECT 3.1125 0.4875 3.1725 0.5475 ;
        RECT 3.0150 0.2475 3.0750 0.3075 ;
        RECT 3.0150 0.7425 3.0750 0.8025 ;
        RECT 2.9100 0.4875 2.9700 0.5475 ;
        RECT 2.8050 0.1200 2.8650 0.1800 ;
        RECT 2.8050 0.8700 2.8650 0.9300 ;
        RECT 2.7000 0.4875 2.7600 0.5475 ;
        RECT 2.5950 0.8100 2.6550 0.8700 ;
        RECT 2.4900 0.4725 2.5500 0.5325 ;
        RECT 2.3850 0.2250 2.4450 0.2850 ;
        RECT 2.3850 0.8325 2.4450 0.8925 ;
        RECT 2.1750 0.2700 2.2350 0.3300 ;
        RECT 2.1750 0.7200 2.2350 0.7800 ;
        RECT 2.0700 0.4725 2.1300 0.5325 ;
        RECT 1.9650 0.1200 2.0250 0.1800 ;
        RECT 1.9650 0.8625 2.0250 0.9225 ;
        RECT 1.8675 0.4650 1.9275 0.5250 ;
        RECT 1.7550 0.2325 1.8150 0.2925 ;
        RECT 1.7550 0.6525 1.8150 0.7125 ;
        RECT 1.5450 0.1575 1.6050 0.2175 ;
        RECT 1.5450 0.8325 1.6050 0.8925 ;
        RECT 1.4325 0.6450 1.4925 0.7050 ;
        RECT 1.3350 0.1275 1.3950 0.1875 ;
        RECT 1.3350 0.8700 1.3950 0.9300 ;
        RECT 1.2300 0.3150 1.2900 0.3750 ;
        RECT 1.0200 0.3525 1.0800 0.4125 ;
        RECT 1.0200 0.6150 1.0800 0.6750 ;
        RECT 0.9150 0.1575 0.9750 0.2175 ;
        RECT 0.9150 0.8325 0.9750 0.8925 ;
        RECT 0.8175 0.3975 0.8775 0.4575 ;
        RECT 0.7050 0.1575 0.7650 0.2175 ;
        RECT 0.7050 0.8100 0.7650 0.8700 ;
        RECT 0.6075 0.5775 0.6675 0.6375 ;
        RECT 0.4950 0.2100 0.5550 0.2700 ;
        RECT 0.4950 0.8100 0.5550 0.8700 ;
        RECT 0.3900 0.4650 0.4500 0.5250 ;
        RECT 0.2850 0.1200 0.3450 0.1800 ;
        RECT 0.1725 0.4650 0.2325 0.5250 ;
        RECT 0.0750 0.2100 0.1350 0.2700 ;
        RECT 0.0750 0.8325 0.1350 0.8925 ;
        LAYER M1 ;
        RECT 2.9325 0.4575 3.1725 0.5775 ;
        RECT 2.8575 0.2550 2.9325 0.7950 ;
        RECT 2.4525 0.2550 2.8575 0.3300 ;
        RECT 2.6775 0.7200 2.8575 0.7950 ;
        RECT 2.6250 0.4050 2.7825 0.6450 ;
        RECT 2.5725 0.7200 2.6775 0.8925 ;
        RECT 2.3925 0.4425 2.5500 0.5625 ;
        RECT 2.3775 0.1800 2.4525 0.3300 ;
        RECT 2.2275 0.4125 2.3925 0.5625 ;
        RECT 1.9950 0.2625 2.2650 0.3375 ;
        RECT 1.9950 0.7125 2.2650 0.7875 ;
        RECT 2.0700 0.4425 2.2275 0.5625 ;
        RECT 1.9200 0.2625 1.9950 0.7875 ;
        RECT 1.8675 0.4350 1.9200 0.5550 ;
        RECT 1.7925 0.2025 1.8375 0.3225 ;
        RECT 1.7925 0.6300 1.8375 0.7350 ;
        RECT 1.7175 0.2025 1.7925 0.7350 ;
        RECT 1.5675 0.1500 1.6425 0.9000 ;
        RECT 1.5150 0.1500 1.5675 0.3600 ;
        RECT 1.5150 0.8250 1.5675 0.9000 ;
        RECT 1.2975 0.2850 1.5150 0.3600 ;
        RECT 1.2600 0.6150 1.4925 0.7350 ;
        RECT 1.2225 0.2850 1.2975 0.4050 ;
        RECT 1.1850 0.6150 1.2600 0.9000 ;
        RECT 0.8850 0.8100 1.1850 0.9000 ;
        RECT 1.0200 0.3225 1.1400 0.4875 ;
        RECT 0.9150 0.5625 1.0800 0.7050 ;
        RECT 0.8175 0.3675 1.0200 0.4875 ;
        RECT 0.7425 0.1500 1.0125 0.2250 ;
        RECT 0.6975 0.6150 0.9150 0.7050 ;
        RECT 0.4875 0.7800 0.7800 0.9000 ;
        RECT 0.6675 0.1500 0.7425 0.5025 ;
        RECT 0.5775 0.5775 0.6975 0.7050 ;
        RECT 0.5775 0.4125 0.6675 0.5025 ;
        RECT 0.4875 0.1800 0.5625 0.3300 ;
        RECT 0.1425 0.2550 0.4875 0.3300 ;
        RECT 0.3075 0.4050 0.4725 0.6000 ;
        RECT 0.2475 0.6750 0.3825 0.8175 ;
        RECT 0.2325 0.6750 0.2475 0.7500 ;
        RECT 0.1575 0.4350 0.2325 0.7500 ;
        RECT 0.0675 0.1800 0.1425 0.3300 ;
        LAYER VIA1 ;
        RECT 2.6775 0.5250 2.7525 0.6000 ;
        RECT 1.9200 0.5625 1.9950 0.6375 ;
        RECT 1.7175 0.3675 1.7925 0.4425 ;
        RECT 1.5675 0.7125 1.6425 0.7875 ;
        RECT 1.1850 0.7125 1.2600 0.7875 ;
        RECT 1.0650 0.3675 1.1400 0.4425 ;
        RECT 0.9600 0.5625 1.0350 0.6375 ;
        RECT 0.6225 0.4275 0.6975 0.5025 ;
        LAYER M2 ;
        RECT 2.6775 0.4800 2.7525 0.7875 ;
        RECT 1.5225 0.7125 2.6775 0.7875 ;
        RECT 0.9150 0.5625 2.0400 0.6375 ;
        RECT 1.0200 0.3675 1.8375 0.4425 ;
        RECT 0.7650 0.7125 1.3050 0.7875 ;
        RECT 0.6900 0.4275 0.7650 0.7875 ;
        RECT 0.5775 0.4275 0.6900 0.5025 ;
    END
END CKLNQ_0011


MACRO CKLNQ_0100
    CLASS CORE ;
    FOREIGN CKLNQ_0100 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.8300 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN TE
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.0900 0.7125 0.5700 0.7875 ;
        VIA 0.3150 0.7500 VIA12_square ;
        END
    END TE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 3.8325 0.2775 3.9900 0.3975 ;
        RECT 3.8325 0.6225 3.9900 0.7425 ;
        RECT 3.5175 0.2775 3.8325 0.7425 ;
        RECT 3.3600 0.2775 3.5175 0.3975 ;
        RECT 3.3600 0.6225 3.5175 0.7425 ;
        VIA 3.8325 0.3375 VIA12_slot ;
        VIA 3.8325 0.6825 VIA12_slot ;
        VIA 3.5175 0.3375 VIA12_slot ;
        VIA 3.5175 0.6825 VIA12_slot ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.4275 0.2625 0.8925 0.3375 ;
        RECT 0.3525 0.2625 0.4275 0.5400 ;
        VIA 0.3900 0.4575 VIA12_square ;
        END
    END E
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 4.2150 0.4125 4.6875 0.4875 ;
        RECT 4.1400 0.1125 4.2150 0.4875 ;
        RECT 2.4825 0.1125 4.1400 0.1875 ;
        RECT 2.3775 0.1125 2.4825 0.5925 ;
        VIA 4.5750 0.4500 VIA12_square ;
        VIA 2.4300 0.5100 VIA12_square ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 4.5600 -0.0750 4.8300 0.0750 ;
        RECT 4.4550 -0.0750 4.5600 0.2400 ;
        RECT 4.1550 -0.0750 4.4550 0.0750 ;
        RECT 4.0350 -0.0750 4.1550 0.2025 ;
        RECT 3.7350 -0.0750 4.0350 0.0750 ;
        RECT 3.6150 -0.0750 3.7350 0.2025 ;
        RECT 3.3150 -0.0750 3.6150 0.0750 ;
        RECT 3.1950 -0.0750 3.3150 0.2025 ;
        RECT 2.8950 -0.0750 3.1950 0.0750 ;
        RECT 2.7900 -0.0750 2.8950 0.2250 ;
        RECT 2.0400 -0.0750 2.7900 0.0750 ;
        RECT 1.9500 -0.0750 2.0400 0.2325 ;
        RECT 1.4250 -0.0750 1.9500 0.0750 ;
        RECT 1.3050 -0.0750 1.4250 0.2100 ;
        RECT 0.3750 -0.0750 1.3050 0.0750 ;
        RECT 0.2550 -0.0750 0.3750 0.1800 ;
        RECT 0.0000 -0.0750 0.2550 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 4.5750 0.9750 4.8300 1.1250 ;
        RECT 4.4550 0.8625 4.5750 1.1250 ;
        RECT 4.1550 0.9750 4.4550 1.1250 ;
        RECT 4.0350 0.8250 4.1550 1.1250 ;
        RECT 3.7350 0.9750 4.0350 1.1250 ;
        RECT 3.6150 0.8250 3.7350 1.1250 ;
        RECT 3.3150 0.9750 3.6150 1.1250 ;
        RECT 3.1950 0.8250 3.3150 1.1250 ;
        RECT 2.8950 0.9750 3.1950 1.1250 ;
        RECT 2.7750 0.8700 2.8950 1.1250 ;
        RECT 2.4750 0.9750 2.7750 1.1250 ;
        RECT 2.3550 0.8700 2.4750 1.1250 ;
        RECT 2.0550 0.9750 2.3550 1.1250 ;
        RECT 1.9350 0.8625 2.0550 1.1250 ;
        RECT 1.4100 0.9750 1.9350 1.1250 ;
        RECT 1.3350 0.8400 1.4100 1.1250 ;
        RECT 0.1650 0.9750 1.3350 1.1250 ;
        RECT 0.0450 0.8250 0.1650 1.1250 ;
        RECT 0.0000 0.9750 0.0450 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 4.6950 0.1725 4.7550 0.2325 ;
        RECT 4.6950 0.7200 4.7550 0.7800 ;
        RECT 4.5825 0.4800 4.6425 0.5400 ;
        RECT 4.4850 0.1500 4.5450 0.2100 ;
        RECT 4.4850 0.8700 4.5450 0.9300 ;
        RECT 4.3725 0.4875 4.4325 0.5475 ;
        RECT 4.2750 0.3075 4.3350 0.3675 ;
        RECT 4.2750 0.7875 4.3350 0.8475 ;
        RECT 4.1700 0.4800 4.2300 0.5400 ;
        RECT 4.0650 0.1350 4.1250 0.1950 ;
        RECT 4.0650 0.8325 4.1250 0.8925 ;
        RECT 3.9600 0.4800 4.0200 0.5400 ;
        RECT 3.8550 0.3075 3.9150 0.3675 ;
        RECT 3.8550 0.6525 3.9150 0.7125 ;
        RECT 3.7500 0.4800 3.8100 0.5400 ;
        RECT 3.6450 0.1350 3.7050 0.1950 ;
        RECT 3.6450 0.8325 3.7050 0.8925 ;
        RECT 3.5400 0.4800 3.6000 0.5400 ;
        RECT 3.4350 0.3075 3.4950 0.3675 ;
        RECT 3.4350 0.6525 3.4950 0.7125 ;
        RECT 3.3300 0.4800 3.3900 0.5400 ;
        RECT 3.2250 0.1350 3.2850 0.1950 ;
        RECT 3.2250 0.8325 3.2850 0.8925 ;
        RECT 3.1200 0.4800 3.1800 0.5400 ;
        RECT 3.0150 0.3075 3.0750 0.3675 ;
        RECT 3.0150 0.6525 3.0750 0.7125 ;
        RECT 2.9100 0.4800 2.9700 0.5400 ;
        RECT 2.8050 0.1350 2.8650 0.1950 ;
        RECT 2.8050 0.8700 2.8650 0.9300 ;
        RECT 2.7000 0.4950 2.7600 0.5550 ;
        RECT 2.5950 0.1575 2.6550 0.2175 ;
        RECT 2.5950 0.8100 2.6550 0.8700 ;
        RECT 2.4900 0.4875 2.5500 0.5475 ;
        RECT 2.3850 0.3075 2.4450 0.3675 ;
        RECT 2.3850 0.8700 2.4450 0.9300 ;
        RECT 2.2800 0.4875 2.3400 0.5475 ;
        RECT 2.1750 0.1575 2.2350 0.2175 ;
        RECT 2.1750 0.8100 2.2350 0.8700 ;
        RECT 2.0700 0.4875 2.1300 0.5475 ;
        RECT 1.9650 0.1425 2.0250 0.2025 ;
        RECT 1.9650 0.8625 2.0250 0.9225 ;
        RECT 1.8675 0.4650 1.9275 0.5250 ;
        RECT 1.7550 0.2325 1.8150 0.2925 ;
        RECT 1.7550 0.6525 1.8150 0.7125 ;
        RECT 1.5450 0.1575 1.6050 0.2175 ;
        RECT 1.5450 0.8325 1.6050 0.8925 ;
        RECT 1.4325 0.6450 1.4925 0.7050 ;
        RECT 1.3350 0.1275 1.3950 0.1875 ;
        RECT 1.3350 0.8700 1.3950 0.9300 ;
        RECT 1.2300 0.3150 1.2900 0.3750 ;
        RECT 1.0200 0.3525 1.0800 0.4125 ;
        RECT 1.0200 0.6150 1.0800 0.6750 ;
        RECT 0.9150 0.1575 0.9750 0.2175 ;
        RECT 0.9150 0.8325 0.9750 0.8925 ;
        RECT 0.8175 0.3975 0.8775 0.4575 ;
        RECT 0.7050 0.1575 0.7650 0.2175 ;
        RECT 0.7050 0.8100 0.7650 0.8700 ;
        RECT 0.6075 0.5775 0.6675 0.6375 ;
        RECT 0.4950 0.2100 0.5550 0.2700 ;
        RECT 0.4950 0.8100 0.5550 0.8700 ;
        RECT 0.3900 0.4650 0.4500 0.5250 ;
        RECT 0.2850 0.1200 0.3450 0.1800 ;
        RECT 0.1725 0.4650 0.2325 0.5250 ;
        RECT 0.0750 0.2100 0.1350 0.2700 ;
        RECT 0.0750 0.8325 0.1350 0.8925 ;
        LAYER M1 ;
        RECT 4.7175 0.1500 4.7925 0.7875 ;
        RECT 4.6650 0.1500 4.7175 0.2400 ;
        RECT 4.4400 0.7125 4.7175 0.7875 ;
        RECT 4.5375 0.3150 4.6425 0.6075 ;
        RECT 4.4400 0.3150 4.5375 0.3975 ;
        RECT 4.3800 0.4725 4.4625 0.5775 ;
        RECT 2.9400 0.4725 4.3800 0.5475 ;
        RECT 3.0150 0.2775 4.3350 0.3975 ;
        RECT 4.3050 0.7575 4.3350 0.8775 ;
        RECT 4.2300 0.6225 4.3050 0.8775 ;
        RECT 3.0150 0.6225 4.2300 0.7425 ;
        RECT 2.8650 0.3000 2.9400 0.7950 ;
        RECT 2.3550 0.3000 2.8650 0.3750 ;
        RECT 2.6775 0.7200 2.8650 0.7950 ;
        RECT 2.6250 0.4500 2.7900 0.6450 ;
        RECT 2.1450 0.1500 2.6850 0.2250 ;
        RECT 2.5725 0.7200 2.6775 0.8925 ;
        RECT 2.2575 0.7200 2.5725 0.7950 ;
        RECT 2.2725 0.4500 2.5500 0.5775 ;
        RECT 2.1525 0.7200 2.2575 0.8925 ;
        RECT 2.0700 0.3450 2.1825 0.6450 ;
        RECT 1.9200 0.3375 1.9950 0.7575 ;
        RECT 1.8675 0.4350 1.9200 0.5550 ;
        RECT 1.7925 0.2025 1.8375 0.3225 ;
        RECT 1.7925 0.6300 1.8375 0.7350 ;
        RECT 1.7175 0.2025 1.7925 0.7350 ;
        RECT 1.5675 0.1500 1.6425 0.9000 ;
        RECT 1.5150 0.1500 1.5675 0.3600 ;
        RECT 1.5150 0.8250 1.5675 0.9000 ;
        RECT 1.2975 0.2850 1.5150 0.3600 ;
        RECT 1.2600 0.6150 1.4925 0.7350 ;
        RECT 1.2225 0.2850 1.2975 0.4050 ;
        RECT 1.1850 0.6150 1.2600 0.9000 ;
        RECT 0.8850 0.8100 1.1850 0.9000 ;
        RECT 1.0200 0.3225 1.1400 0.4875 ;
        RECT 0.9150 0.5625 1.0800 0.7050 ;
        RECT 0.8175 0.3675 1.0200 0.4875 ;
        RECT 0.7425 0.1500 1.0125 0.2250 ;
        RECT 0.6975 0.6150 0.9150 0.7050 ;
        RECT 0.4875 0.7800 0.7800 0.9000 ;
        RECT 0.6675 0.1500 0.7425 0.5025 ;
        RECT 0.5775 0.5775 0.6975 0.7050 ;
        RECT 0.5775 0.4125 0.6675 0.5025 ;
        RECT 0.4875 0.1800 0.5625 0.3300 ;
        RECT 0.1425 0.2550 0.4875 0.3300 ;
        RECT 0.3075 0.4050 0.4725 0.6000 ;
        RECT 0.2475 0.6750 0.3825 0.8175 ;
        RECT 0.2325 0.6750 0.2475 0.7500 ;
        RECT 0.1575 0.4350 0.2325 0.7500 ;
        RECT 0.0675 0.1800 0.1425 0.3300 ;
        LAYER VIA1 ;
        RECT 4.4850 0.7125 4.5600 0.7875 ;
        RECT 2.6775 0.4950 2.7525 0.5700 ;
        RECT 2.1075 0.4125 2.1825 0.4875 ;
        RECT 1.9200 0.6225 1.9950 0.6975 ;
        RECT 1.7175 0.4125 1.7925 0.4875 ;
        RECT 1.5675 0.2625 1.6425 0.3375 ;
        RECT 1.1850 0.7125 1.2600 0.7875 ;
        RECT 1.0650 0.3675 1.1400 0.4425 ;
        RECT 0.9600 0.5625 1.0350 0.6375 ;
        RECT 0.6225 0.4275 0.6975 0.5025 ;
        LAYER M2 ;
        RECT 3.8625 0.2775 3.9900 0.3975 ;
        RECT 3.8625 0.6225 3.9900 0.7425 ;
        RECT 3.3600 0.2775 3.4875 0.3975 ;
        RECT 3.3600 0.6225 3.4875 0.7425 ;
        RECT 4.2150 0.7125 4.6350 0.7875 ;
        RECT 4.1400 0.7125 4.2150 0.9375 ;
        RECT 1.9950 0.8625 4.1400 0.9375 ;
        RECT 2.6775 0.4500 2.7525 0.7875 ;
        RECT 2.1825 0.7125 2.6775 0.7875 ;
        RECT 2.1075 0.2625 2.1825 0.7875 ;
        RECT 1.4925 0.2625 2.1075 0.3375 ;
        RECT 1.9200 0.5625 1.9950 0.9375 ;
        RECT 0.9150 0.5625 1.9200 0.6375 ;
        RECT 1.3425 0.4125 1.8675 0.4875 ;
        RECT 1.2600 0.3675 1.3425 0.4875 ;
        RECT 0.7650 0.7125 1.3050 0.7875 ;
        RECT 1.0200 0.3675 1.2600 0.4425 ;
        RECT 0.6900 0.4275 0.7650 0.7875 ;
        RECT 0.5775 0.4275 0.6900 0.5025 ;
    END
END CKLNQ_0100


MACRO CKLNQ_0101
    CLASS CORE ;
    FOREIGN CKLNQ_0101 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.9300 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN TE
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.9975 0.2625 1.0725 0.6450 ;
        RECT 0.3225 0.2625 0.9975 0.3375 ;
        VIA 1.0350 0.5625 VIA12_square ;
        VIA 0.4575 0.3000 VIA12_square ;
        END
    END TE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 5.0850 0.2775 5.2425 0.3975 ;
        RECT 5.0850 0.6300 5.2425 0.7500 ;
        RECT 4.7700 0.2775 5.0850 0.7500 ;
        RECT 4.6125 0.2775 4.7700 0.3975 ;
        RECT 4.6125 0.6300 4.7700 0.7500 ;
        VIA 5.0850 0.3375 VIA12_slot ;
        VIA 5.0850 0.6900 VIA12_slot ;
        VIA 4.7700 0.3375 VIA12_slot ;
        VIA 4.7700 0.6900 VIA12_slot ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.2075 0.1125 1.3125 0.6225 ;
        RECT 0.7575 0.1125 1.2075 0.1875 ;
        VIA 1.2600 0.5325 VIA12_square ;
        END
    END E
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 6.1500 0.4125 6.6525 0.4875 ;
        RECT 6.0450 0.4125 6.1500 0.6075 ;
        VIA 6.0975 0.5250 VIA12_square ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 5.8275 -0.0750 6.9300 0.0750 ;
        RECT 5.7225 -0.0750 5.8275 0.2100 ;
        RECT 5.4150 -0.0750 5.7225 0.0750 ;
        RECT 5.2950 -0.0750 5.4150 0.1800 ;
        RECT 4.9950 -0.0750 5.2950 0.0750 ;
        RECT 4.8750 -0.0750 4.9950 0.1800 ;
        RECT 4.5750 -0.0750 4.8750 0.0750 ;
        RECT 4.4550 -0.0750 4.5750 0.1800 ;
        RECT 4.1550 -0.0750 4.4550 0.0750 ;
        RECT 4.0350 -0.0750 4.1550 0.1800 ;
        RECT 3.7350 -0.0750 4.0350 0.0750 ;
        RECT 3.6150 -0.0750 3.7350 0.1800 ;
        RECT 3.3150 -0.0750 3.6150 0.0750 ;
        RECT 3.1950 -0.0750 3.3150 0.1800 ;
        RECT 2.7000 -0.0750 3.1950 0.0750 ;
        RECT 2.5950 -0.0750 2.7000 0.2625 ;
        RECT 1.8150 -0.0750 2.5950 0.0750 ;
        RECT 1.7100 -0.0750 1.8150 0.2250 ;
        RECT 0.3450 -0.0750 1.7100 0.0750 ;
        RECT 0.2400 -0.0750 0.3450 0.2250 ;
        RECT 0.0000 -0.0750 0.2400 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 6.8775 0.9750 6.9300 1.1250 ;
        RECT 6.7725 0.8100 6.8775 1.1250 ;
        RECT 6.4800 0.9750 6.7725 1.1250 ;
        RECT 6.3750 0.8100 6.4800 1.1250 ;
        RECT 5.8050 0.9750 6.3750 1.1250 ;
        RECT 5.7000 0.8100 5.8050 1.1250 ;
        RECT 5.4150 0.9750 5.7000 1.1250 ;
        RECT 5.2950 0.8250 5.4150 1.1250 ;
        RECT 4.9950 0.9750 5.2950 1.1250 ;
        RECT 4.8750 0.8250 4.9950 1.1250 ;
        RECT 4.5750 0.9750 4.8750 1.1250 ;
        RECT 4.4550 0.8250 4.5750 1.1250 ;
        RECT 4.1550 0.9750 4.4550 1.1250 ;
        RECT 4.0350 0.8250 4.1550 1.1250 ;
        RECT 3.7350 0.9750 4.0350 1.1250 ;
        RECT 3.6150 0.8250 3.7350 1.1250 ;
        RECT 3.3150 0.9750 3.6150 1.1250 ;
        RECT 3.1950 0.8250 3.3150 1.1250 ;
        RECT 2.8950 0.9750 3.1950 1.1250 ;
        RECT 2.7750 0.8325 2.8950 1.1250 ;
        RECT 2.0550 0.9750 2.7750 1.1250 ;
        RECT 1.9350 0.8250 2.0550 1.1250 ;
        RECT 0.7950 0.9750 1.9350 1.1250 ;
        RECT 0.6750 0.8625 0.7950 1.1250 ;
        RECT 0.3600 0.9750 0.6750 1.1250 ;
        RECT 0.2550 0.8250 0.3600 1.1250 ;
        RECT 0.0000 0.9750 0.2550 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 6.7950 0.3075 6.8550 0.3675 ;
        RECT 6.7950 0.8325 6.8550 0.8925 ;
        RECT 6.6825 0.4950 6.7425 0.5550 ;
        RECT 6.5850 0.1650 6.6450 0.2250 ;
        RECT 6.5850 0.8100 6.6450 0.8700 ;
        RECT 6.4800 0.4950 6.5400 0.5550 ;
        RECT 6.3750 0.3075 6.4350 0.3675 ;
        RECT 6.3750 0.8475 6.4350 0.9075 ;
        RECT 6.2700 0.4950 6.3300 0.5550 ;
        RECT 6.1650 0.1650 6.2250 0.2250 ;
        RECT 6.1650 0.6750 6.2250 0.7350 ;
        RECT 5.9550 0.2475 6.0150 0.3075 ;
        RECT 5.9550 0.8250 6.0150 0.8850 ;
        RECT 5.8500 0.4950 5.9100 0.5550 ;
        RECT 5.7450 0.1200 5.8050 0.1800 ;
        RECT 5.7450 0.8475 5.8050 0.9075 ;
        RECT 5.6400 0.4800 5.7000 0.5400 ;
        RECT 5.5350 0.3000 5.5950 0.3600 ;
        RECT 5.5350 0.6600 5.5950 0.7200 ;
        RECT 5.4300 0.4800 5.4900 0.5400 ;
        RECT 5.3250 0.1200 5.3850 0.1800 ;
        RECT 5.3250 0.8325 5.3850 0.8925 ;
        RECT 5.2200 0.4800 5.2800 0.5400 ;
        RECT 5.1150 0.3000 5.1750 0.3600 ;
        RECT 5.1150 0.6600 5.1750 0.7200 ;
        RECT 5.0100 0.4800 5.0700 0.5400 ;
        RECT 4.9050 0.1200 4.9650 0.1800 ;
        RECT 4.9050 0.8325 4.9650 0.8925 ;
        RECT 4.8000 0.4800 4.8600 0.5400 ;
        RECT 4.6950 0.3000 4.7550 0.3600 ;
        RECT 4.6950 0.6600 4.7550 0.7200 ;
        RECT 4.5900 0.4800 4.6500 0.5400 ;
        RECT 4.4850 0.1200 4.5450 0.1800 ;
        RECT 4.4850 0.8325 4.5450 0.8925 ;
        RECT 4.3800 0.4800 4.4400 0.5400 ;
        RECT 4.2750 0.3000 4.3350 0.3600 ;
        RECT 4.2750 0.6600 4.3350 0.7200 ;
        RECT 4.1700 0.4800 4.2300 0.5400 ;
        RECT 4.0650 0.1200 4.1250 0.1800 ;
        RECT 4.0650 0.8325 4.1250 0.8925 ;
        RECT 3.9600 0.4950 4.0200 0.5550 ;
        RECT 3.8550 0.2700 3.9150 0.3300 ;
        RECT 3.8550 0.6750 3.9150 0.7350 ;
        RECT 3.7500 0.4950 3.8100 0.5550 ;
        RECT 3.6450 0.1200 3.7050 0.1800 ;
        RECT 3.6450 0.8325 3.7050 0.8925 ;
        RECT 3.5400 0.4950 3.6000 0.5550 ;
        RECT 3.4350 0.2700 3.4950 0.3300 ;
        RECT 3.3300 0.4950 3.3900 0.5550 ;
        RECT 3.2250 0.1200 3.2850 0.1800 ;
        RECT 3.2250 0.8325 3.2850 0.8925 ;
        RECT 3.1275 0.4875 3.1875 0.5475 ;
        RECT 3.0150 0.2550 3.0750 0.3150 ;
        RECT 3.0150 0.7500 3.0750 0.8100 ;
        RECT 2.8050 0.1725 2.8650 0.2325 ;
        RECT 2.8050 0.8325 2.8650 0.8925 ;
        RECT 2.6925 0.4650 2.7525 0.5250 ;
        RECT 2.5950 0.1725 2.6550 0.2325 ;
        RECT 2.5950 0.6900 2.6550 0.7500 ;
        RECT 2.4900 0.4650 2.5500 0.5250 ;
        RECT 2.3850 0.1725 2.4450 0.2325 ;
        RECT 2.1750 0.1800 2.2350 0.2400 ;
        RECT 2.1750 0.8325 2.2350 0.8925 ;
        RECT 2.0700 0.3675 2.1300 0.4275 ;
        RECT 1.9650 0.8325 2.0250 0.8925 ;
        RECT 1.8600 0.5250 1.9200 0.5850 ;
        RECT 1.7550 0.1275 1.8150 0.1875 ;
        RECT 1.6500 0.5550 1.7100 0.6150 ;
        RECT 1.5450 0.1725 1.6050 0.2325 ;
        RECT 1.5450 0.8325 1.6050 0.8925 ;
        RECT 1.3350 0.1575 1.3950 0.2175 ;
        RECT 1.3350 0.8175 1.3950 0.8775 ;
        RECT 1.2300 0.4800 1.2900 0.5400 ;
        RECT 1.1250 0.3000 1.1850 0.3600 ;
        RECT 1.1250 0.8175 1.1850 0.8775 ;
        RECT 1.0200 0.4800 1.0800 0.5400 ;
        RECT 0.9150 0.1950 0.9750 0.2550 ;
        RECT 0.9150 0.8100 0.9750 0.8700 ;
        RECT 0.8100 0.4875 0.8700 0.5475 ;
        RECT 0.7050 0.1725 0.7650 0.2325 ;
        RECT 0.7050 0.8700 0.7650 0.9300 ;
        RECT 0.6000 0.4950 0.6600 0.5550 ;
        RECT 0.4950 0.8325 0.5550 0.8925 ;
        RECT 0.3900 0.4875 0.4500 0.5475 ;
        RECT 0.2850 0.1350 0.3450 0.1950 ;
        RECT 0.2850 0.8550 0.3450 0.9150 ;
        RECT 0.1875 0.4800 0.2475 0.5400 ;
        RECT 0.0750 0.2625 0.1350 0.3225 ;
        RECT 0.0750 0.6900 0.1350 0.7500 ;
        LAYER M1 ;
        RECT 6.8175 0.3075 6.8925 0.7350 ;
        RECT 6.3375 0.3075 6.8175 0.3900 ;
        RECT 6.6675 0.6600 6.8175 0.7350 ;
        RECT 6.3225 0.4650 6.7425 0.5850 ;
        RECT 6.1275 0.1575 6.6900 0.2325 ;
        RECT 6.5625 0.6600 6.6675 0.9000 ;
        RECT 5.7525 0.6600 6.5625 0.7350 ;
        RECT 5.8275 0.4725 6.3225 0.5850 ;
        RECT 5.9100 0.8100 6.2700 0.9000 ;
        RECT 5.9475 0.1950 6.0225 0.3975 ;
        RECT 5.7225 0.3000 5.9475 0.3975 ;
        RECT 5.6775 0.4800 5.7525 0.7350 ;
        RECT 4.1775 0.4800 5.6775 0.5550 ;
        RECT 4.2450 0.2775 5.6175 0.3975 ;
        RECT 4.2675 0.6300 5.5950 0.7500 ;
        RECT 4.1025 0.4800 4.1775 0.7425 ;
        RECT 3.3225 0.2550 4.1250 0.3750 ;
        RECT 3.7875 0.6675 4.1025 0.7425 ;
        RECT 3.3225 0.4650 4.0275 0.5850 ;
        RECT 3.1575 0.4200 3.2475 0.7200 ;
        RECT 3.1275 0.4200 3.1575 0.6225 ;
        RECT 3.0525 0.2250 3.0975 0.3375 ;
        RECT 3.0525 0.7200 3.0825 0.8400 ;
        RECT 2.9775 0.2250 3.0525 0.8400 ;
        RECT 2.8275 0.1500 2.9025 0.7575 ;
        RECT 2.7825 0.1500 2.8275 0.2550 ;
        RECT 2.4075 0.6825 2.8275 0.7575 ;
        RECT 2.6325 0.3450 2.7525 0.6075 ;
        RECT 2.4825 0.3750 2.5575 0.5775 ;
        RECT 2.3100 0.1500 2.5200 0.3000 ;
        RECT 2.1525 0.3750 2.4825 0.4500 ;
        RECT 2.3325 0.5250 2.4075 0.7575 ;
        RECT 1.8225 0.5250 2.3325 0.6000 ;
        RECT 2.2125 0.8250 2.2650 0.9000 ;
        RECT 1.9650 0.1500 2.2350 0.2700 ;
        RECT 2.1375 0.6750 2.2125 0.9000 ;
        RECT 2.0400 0.3450 2.1525 0.4500 ;
        RECT 1.7100 0.6750 2.1375 0.7500 ;
        RECT 1.8900 0.1500 1.9650 0.4050 ;
        RECT 1.4550 0.3300 1.8900 0.4050 ;
        RECT 1.6350 0.5025 1.7100 0.7500 ;
        RECT 1.4550 0.8250 1.6500 0.9000 ;
        RECT 1.5225 0.1500 1.6275 0.2550 ;
        RECT 0.9825 0.1500 1.5225 0.2250 ;
        RECT 1.3800 0.3000 1.4550 0.9000 ;
        RECT 1.0875 0.3000 1.3800 0.3750 ;
        RECT 1.3125 0.7950 1.3800 0.9000 ;
        RECT 1.1850 0.4500 1.3050 0.7200 ;
        RECT 1.0125 0.7950 1.2075 0.9000 ;
        RECT 0.9525 0.4500 1.1100 0.6975 ;
        RECT 0.9075 0.7725 1.0125 0.9000 ;
        RECT 0.9075 0.1500 0.9825 0.3150 ;
        RECT 0.8250 0.4575 0.8775 0.5850 ;
        RECT 0.7500 0.1500 0.8250 0.7875 ;
        RECT 0.6825 0.1500 0.7500 0.2550 ;
        RECT 0.6000 0.7125 0.7500 0.7875 ;
        RECT 0.5700 0.3375 0.6750 0.6375 ;
        RECT 0.5250 0.7125 0.6000 0.9000 ;
        RECT 0.4650 0.8250 0.5250 0.9000 ;
        RECT 0.4200 0.1950 0.4950 0.3825 ;
        RECT 0.4425 0.4575 0.4725 0.5775 ;
        RECT 0.3675 0.4575 0.4425 0.7500 ;
        RECT 0.2925 0.3075 0.4200 0.3825 ;
        RECT 0.1125 0.6750 0.3675 0.7500 ;
        RECT 0.2175 0.3075 0.2925 0.5700 ;
        RECT 0.1875 0.4350 0.2175 0.5700 ;
        RECT 0.1125 0.2100 0.1425 0.3525 ;
        RECT 0.0375 0.2100 0.1125 0.7500 ;
        LAYER VIA1 ;
        RECT 6.1725 0.1575 6.2475 0.2325 ;
        RECT 5.9550 0.8175 6.0300 0.8925 ;
        RECT 5.7825 0.3225 5.8575 0.3975 ;
        RECT 3.9900 0.2700 4.0650 0.3450 ;
        RECT 3.3825 0.5025 3.4575 0.5775 ;
        RECT 3.1575 0.6000 3.2325 0.6750 ;
        RECT 2.9775 0.3450 3.0525 0.4200 ;
        RECT 2.8275 0.1950 2.9025 0.2700 ;
        RECT 2.6625 0.4950 2.7375 0.5700 ;
        RECT 2.3775 0.1575 2.4525 0.2325 ;
        RECT 2.3625 0.3750 2.4375 0.4500 ;
        RECT 1.6350 0.5625 1.7100 0.6375 ;
        RECT 1.3800 0.7125 1.4550 0.7875 ;
        RECT 0.5775 0.4650 0.6525 0.5400 ;
        LAYER M2 ;
        RECT 5.1150 0.2775 5.2425 0.3975 ;
        RECT 5.1150 0.6300 5.2425 0.7500 ;
        RECT 4.6125 0.2775 4.7400 0.3975 ;
        RECT 4.6125 0.6300 4.7400 0.7500 ;
        RECT 5.9100 0.1575 6.2925 0.2325 ;
        RECT 5.9475 0.8175 6.0750 0.9375 ;
        RECT 5.8725 0.3225 5.9475 0.9375 ;
        RECT 5.8350 0.1125 5.9100 0.2325 ;
        RECT 5.7300 0.3225 5.8725 0.3975 ;
        RECT 3.2475 0.8475 5.8725 0.9375 ;
        RECT 4.0875 0.1125 5.8350 0.1875 ;
        RECT 3.9675 0.1125 4.0875 0.4050 ;
        RECT 3.3825 0.1950 3.4575 0.6375 ;
        RECT 2.7600 0.1950 3.3825 0.2700 ;
        RECT 3.1425 0.5550 3.2475 0.9375 ;
        RECT 0.7725 0.8625 3.1425 0.9375 ;
        RECT 2.4825 0.3450 3.1275 0.4200 ;
        RECT 2.6775 0.4950 2.8050 0.5700 ;
        RECT 2.6025 0.4950 2.6775 0.7875 ;
        RECT 1.3275 0.7125 2.6025 0.7875 ;
        RECT 2.1075 0.1575 2.5275 0.2325 ;
        RECT 2.3175 0.3450 2.4825 0.4650 ;
        RECT 2.0325 0.1575 2.1075 0.6375 ;
        RECT 1.5900 0.5625 2.0325 0.6375 ;
        RECT 0.6975 0.4650 0.7725 0.9375 ;
        RECT 0.5025 0.4650 0.6975 0.5400 ;
    END
END CKLNQ_0101


MACRO CKLNQ_0110
    CLASS CORE ;
    FOREIGN CKLNQ_0110 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.6200 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN TE
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.0900 0.7125 0.5700 0.7875 ;
        VIA 0.3150 0.7500 VIA12_square ;
        END
    END TE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 4.0425 0.2775 4.2000 0.3975 ;
        RECT 4.0425 0.6225 4.2000 0.7425 ;
        RECT 3.7275 0.2775 4.0425 0.7425 ;
        RECT 3.5700 0.2775 3.7275 0.3975 ;
        RECT 3.5700 0.6225 3.7275 0.7425 ;
        VIA 4.0425 0.3375 VIA12_slot ;
        VIA 4.0425 0.6825 VIA12_slot ;
        VIA 3.7275 0.3375 VIA12_slot ;
        VIA 3.7275 0.6825 VIA12_slot ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.4275 0.2625 0.8925 0.3375 ;
        RECT 0.3525 0.2625 0.4275 0.5400 ;
        VIA 0.3900 0.4575 VIA12_square ;
        END
    END E
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 2.7825 0.2625 2.8875 0.5925 ;
        RECT 2.3175 0.2625 2.7825 0.3375 ;
        RECT 2.2125 0.2625 2.3175 0.5625 ;
        VIA 2.8350 0.5100 VIA12_square ;
        VIA 2.2650 0.4800 VIA12_square ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 4.5525 -0.0750 4.6200 0.0750 ;
        RECT 4.4775 -0.0750 4.5525 0.3075 ;
        RECT 4.1550 -0.0750 4.4775 0.0750 ;
        RECT 4.0350 -0.0750 4.1550 0.2025 ;
        RECT 3.7350 -0.0750 4.0350 0.0750 ;
        RECT 3.6150 -0.0750 3.7350 0.2025 ;
        RECT 3.3150 -0.0750 3.6150 0.0750 ;
        RECT 3.2100 -0.0750 3.3150 0.2250 ;
        RECT 2.4525 -0.0750 3.2100 0.0750 ;
        RECT 2.3775 -0.0750 2.4525 0.2625 ;
        RECT 2.0550 -0.0750 2.3775 0.0750 ;
        RECT 1.9350 -0.0750 2.0550 0.1875 ;
        RECT 1.4250 -0.0750 1.9350 0.0750 ;
        RECT 1.3050 -0.0750 1.4250 0.2100 ;
        RECT 0.3750 -0.0750 1.3050 0.0750 ;
        RECT 0.2550 -0.0750 0.3750 0.1800 ;
        RECT 0.0000 -0.0750 0.2550 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 4.5675 0.9750 4.6200 1.1250 ;
        RECT 4.4625 0.6375 4.5675 1.1250 ;
        RECT 4.1550 0.9750 4.4625 1.1250 ;
        RECT 4.0350 0.8250 4.1550 1.1250 ;
        RECT 3.7350 0.9750 4.0350 1.1250 ;
        RECT 3.6150 0.8250 3.7350 1.1250 ;
        RECT 3.3150 0.9750 3.6150 1.1250 ;
        RECT 3.1950 0.8700 3.3150 1.1250 ;
        RECT 2.8950 0.9750 3.1950 1.1250 ;
        RECT 2.7750 0.8700 2.8950 1.1250 ;
        RECT 2.4525 0.9750 2.7750 1.1250 ;
        RECT 2.3775 0.7875 2.4525 1.1250 ;
        RECT 2.0550 0.9750 2.3775 1.1250 ;
        RECT 1.9350 0.8625 2.0550 1.1250 ;
        RECT 1.4100 0.9750 1.9350 1.1250 ;
        RECT 1.3350 0.8400 1.4100 1.1250 ;
        RECT 0.1650 0.9750 1.3350 1.1250 ;
        RECT 0.0450 0.8250 0.1650 1.1250 ;
        RECT 0.0000 0.9750 0.0450 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 4.4850 0.2175 4.5450 0.2775 ;
        RECT 4.4850 0.6675 4.5450 0.7275 ;
        RECT 4.4850 0.8325 4.5450 0.8925 ;
        RECT 4.3800 0.4800 4.4400 0.5400 ;
        RECT 4.2750 0.3075 4.3350 0.3675 ;
        RECT 4.2750 0.6525 4.3350 0.7125 ;
        RECT 4.1700 0.4800 4.2300 0.5400 ;
        RECT 4.0650 0.1350 4.1250 0.1950 ;
        RECT 4.0650 0.8325 4.1250 0.8925 ;
        RECT 3.9600 0.4800 4.0200 0.5400 ;
        RECT 3.8550 0.3075 3.9150 0.3675 ;
        RECT 3.8550 0.6525 3.9150 0.7125 ;
        RECT 3.7500 0.4800 3.8100 0.5400 ;
        RECT 3.6450 0.1350 3.7050 0.1950 ;
        RECT 3.6450 0.8325 3.7050 0.8925 ;
        RECT 3.5400 0.4800 3.6000 0.5400 ;
        RECT 3.4350 0.3075 3.4950 0.3675 ;
        RECT 3.4350 0.6525 3.4950 0.7125 ;
        RECT 3.3300 0.4800 3.3900 0.5400 ;
        RECT 3.2250 0.1350 3.2850 0.1950 ;
        RECT 3.2250 0.8700 3.2850 0.9300 ;
        RECT 3.1200 0.4950 3.1800 0.5550 ;
        RECT 3.0150 0.1575 3.0750 0.2175 ;
        RECT 3.0150 0.7950 3.0750 0.8550 ;
        RECT 2.9100 0.4875 2.9700 0.5475 ;
        RECT 2.8050 0.3075 2.8650 0.3675 ;
        RECT 2.8050 0.8700 2.8650 0.9300 ;
        RECT 2.7000 0.4875 2.7600 0.5475 ;
        RECT 2.5950 0.1575 2.6550 0.2175 ;
        RECT 2.5950 0.7950 2.6550 0.8550 ;
        RECT 2.4900 0.4875 2.5500 0.5475 ;
        RECT 2.3850 0.1725 2.4450 0.2325 ;
        RECT 2.3850 0.8325 2.4450 0.8925 ;
        RECT 2.1750 0.2700 2.2350 0.3300 ;
        RECT 2.1750 0.7200 2.2350 0.7800 ;
        RECT 2.0700 0.4725 2.1300 0.5325 ;
        RECT 1.9650 0.1200 2.0250 0.1800 ;
        RECT 1.9650 0.8625 2.0250 0.9225 ;
        RECT 1.8675 0.4650 1.9275 0.5250 ;
        RECT 1.7550 0.2325 1.8150 0.2925 ;
        RECT 1.7550 0.6525 1.8150 0.7125 ;
        RECT 1.5450 0.1575 1.6050 0.2175 ;
        RECT 1.5450 0.8325 1.6050 0.8925 ;
        RECT 1.4325 0.6450 1.4925 0.7050 ;
        RECT 1.3350 0.1275 1.3950 0.1875 ;
        RECT 1.3350 0.8700 1.3950 0.9300 ;
        RECT 1.2300 0.3150 1.2900 0.3750 ;
        RECT 1.0200 0.3525 1.0800 0.4125 ;
        RECT 1.0200 0.6150 1.0800 0.6750 ;
        RECT 0.9150 0.1575 0.9750 0.2175 ;
        RECT 0.9150 0.8325 0.9750 0.8925 ;
        RECT 0.8175 0.3975 0.8775 0.4575 ;
        RECT 0.7050 0.1575 0.7650 0.2175 ;
        RECT 0.7050 0.8100 0.7650 0.8700 ;
        RECT 0.6075 0.5775 0.6675 0.6375 ;
        RECT 0.4950 0.2100 0.5550 0.2700 ;
        RECT 0.4950 0.8100 0.5550 0.8700 ;
        RECT 0.3900 0.4650 0.4500 0.5250 ;
        RECT 0.2850 0.1200 0.3450 0.1800 ;
        RECT 0.1725 0.4650 0.2325 0.5250 ;
        RECT 0.0750 0.2100 0.1350 0.2700 ;
        RECT 0.0750 0.8325 0.1350 0.8925 ;
        LAYER M1 ;
        RECT 3.3600 0.4725 4.4850 0.5475 ;
        RECT 3.4350 0.2775 4.3650 0.3975 ;
        RECT 3.4350 0.6225 4.3650 0.7425 ;
        RECT 3.2850 0.3000 3.3600 0.7950 ;
        RECT 2.7750 0.3000 3.2850 0.3750 ;
        RECT 3.1050 0.7200 3.2850 0.7950 ;
        RECT 3.0450 0.4500 3.2100 0.6450 ;
        RECT 2.5650 0.1500 3.1050 0.2250 ;
        RECT 2.9850 0.7200 3.1050 0.8700 ;
        RECT 2.6850 0.7200 2.9850 0.7950 ;
        RECT 2.6925 0.4500 2.9700 0.5775 ;
        RECT 2.5650 0.7200 2.6850 0.8700 ;
        RECT 2.4375 0.4425 2.6100 0.6450 ;
        RECT 2.0700 0.4425 2.3475 0.5625 ;
        RECT 1.9950 0.2625 2.2650 0.3375 ;
        RECT 1.9950 0.7125 2.2650 0.7875 ;
        RECT 1.9200 0.2625 1.9950 0.7875 ;
        RECT 1.8675 0.4350 1.9200 0.5550 ;
        RECT 1.7925 0.2025 1.8375 0.3225 ;
        RECT 1.7925 0.6300 1.8375 0.7350 ;
        RECT 1.7175 0.2025 1.7925 0.7350 ;
        RECT 1.5675 0.1500 1.6425 0.9000 ;
        RECT 1.5150 0.1500 1.5675 0.3600 ;
        RECT 1.5150 0.8250 1.5675 0.9000 ;
        RECT 1.2975 0.2850 1.5150 0.3600 ;
        RECT 1.2600 0.6150 1.4925 0.7350 ;
        RECT 1.2225 0.2850 1.2975 0.4050 ;
        RECT 1.1850 0.6150 1.2600 0.9000 ;
        RECT 0.8850 0.8100 1.1850 0.9000 ;
        RECT 1.0200 0.3225 1.1400 0.4875 ;
        RECT 0.9150 0.5625 1.0800 0.7050 ;
        RECT 0.8175 0.3675 1.0200 0.4875 ;
        RECT 0.7425 0.1500 1.0125 0.2250 ;
        RECT 0.6975 0.6150 0.9150 0.7050 ;
        RECT 0.4875 0.7800 0.7800 0.9000 ;
        RECT 0.6675 0.1500 0.7425 0.5025 ;
        RECT 0.5775 0.5775 0.6975 0.7050 ;
        RECT 0.5775 0.4125 0.6675 0.5025 ;
        RECT 0.4875 0.1800 0.5625 0.3300 ;
        RECT 0.1425 0.2550 0.4875 0.3300 ;
        RECT 0.3075 0.4050 0.4725 0.6000 ;
        RECT 0.2475 0.6750 0.3825 0.8175 ;
        RECT 0.2325 0.6750 0.2475 0.7500 ;
        RECT 0.1575 0.4350 0.2325 0.7500 ;
        RECT 0.0675 0.1800 0.1425 0.3300 ;
        LAYER VIA1 ;
        RECT 3.0975 0.4950 3.1725 0.5700 ;
        RECT 2.4825 0.5250 2.5575 0.6000 ;
        RECT 1.9200 0.5625 1.9950 0.6375 ;
        RECT 1.7175 0.3675 1.7925 0.4425 ;
        RECT 1.5675 0.7125 1.6425 0.7875 ;
        RECT 1.1850 0.7125 1.2600 0.7875 ;
        RECT 1.0650 0.3675 1.1400 0.4425 ;
        RECT 0.9600 0.5625 1.0350 0.6375 ;
        RECT 0.6225 0.4275 0.6975 0.5025 ;
        LAYER M2 ;
        RECT 4.0725 0.2775 4.2000 0.3975 ;
        RECT 4.0725 0.6225 4.2000 0.7425 ;
        RECT 3.5700 0.2775 3.6975 0.3975 ;
        RECT 3.5700 0.6225 3.6975 0.7425 ;
        RECT 3.0975 0.4500 3.1725 0.7875 ;
        RECT 2.5575 0.7125 3.0975 0.7875 ;
        RECT 2.4825 0.4800 2.5575 0.7875 ;
        RECT 1.5225 0.7125 2.4825 0.7875 ;
        RECT 0.9150 0.5625 2.0400 0.6375 ;
        RECT 1.0200 0.3675 1.8375 0.4425 ;
        RECT 0.7650 0.7125 1.3050 0.7875 ;
        RECT 0.6900 0.4275 0.7650 0.7875 ;
        RECT 0.5775 0.4275 0.6900 0.5025 ;
    END
END CKLNQ_0110


MACRO CKLNQ_0111
    CLASS CORE ;
    FOREIGN CKLNQ_0111 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.7800 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN TE
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.0900 0.7125 0.5700 0.7875 ;
        VIA 0.3150 0.7500 VIA12_square ;
        END
    END TE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 3.0975 0.2550 3.4125 0.7650 ;
        VIA 3.2550 0.3375 VIA12_slot ;
        VIA 3.2550 0.6825 VIA12_slot ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.4275 0.2625 0.8925 0.3375 ;
        RECT 0.3525 0.2625 0.4275 0.5400 ;
        VIA 0.3900 0.4575 VIA12_square ;
        END
    END E
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 2.0250 0.4125 2.4900 0.4875 ;
        VIA 2.3100 0.4500 VIA12_square ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 3.7125 -0.0750 3.7800 0.0750 ;
        RECT 3.6375 -0.0750 3.7125 0.2925 ;
        RECT 3.3150 -0.0750 3.6375 0.0750 ;
        RECT 3.1950 -0.0750 3.3150 0.2025 ;
        RECT 2.8950 -0.0750 3.1950 0.0750 ;
        RECT 2.7750 -0.0750 2.8950 0.1800 ;
        RECT 2.0550 -0.0750 2.7750 0.0750 ;
        RECT 1.9350 -0.0750 2.0550 0.1875 ;
        RECT 1.4250 -0.0750 1.9350 0.0750 ;
        RECT 1.3050 -0.0750 1.4250 0.2100 ;
        RECT 0.3750 -0.0750 1.3050 0.0750 ;
        RECT 0.2550 -0.0750 0.3750 0.1800 ;
        RECT 0.0000 -0.0750 0.2550 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 3.7275 0.9750 3.7800 1.1250 ;
        RECT 3.6225 0.6375 3.7275 1.1250 ;
        RECT 3.3150 0.9750 3.6225 1.1250 ;
        RECT 3.1950 0.8250 3.3150 1.1250 ;
        RECT 2.8950 0.9750 3.1950 1.1250 ;
        RECT 2.7750 0.8700 2.8950 1.1250 ;
        RECT 2.4525 0.9750 2.7750 1.1250 ;
        RECT 2.3775 0.8025 2.4525 1.1250 ;
        RECT 2.0550 0.9750 2.3775 1.1250 ;
        RECT 1.9350 0.8625 2.0550 1.1250 ;
        RECT 1.4100 0.9750 1.9350 1.1250 ;
        RECT 1.3350 0.8400 1.4100 1.1250 ;
        RECT 0.1650 0.9750 1.3350 1.1250 ;
        RECT 0.0450 0.8250 0.1650 1.1250 ;
        RECT 0.0000 0.9750 0.0450 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 3.6450 0.2025 3.7050 0.2625 ;
        RECT 3.6450 0.6675 3.7050 0.7275 ;
        RECT 3.6450 0.8325 3.7050 0.8925 ;
        RECT 3.5400 0.4800 3.6000 0.5400 ;
        RECT 3.4350 0.3075 3.4950 0.3675 ;
        RECT 3.4350 0.6525 3.4950 0.7125 ;
        RECT 3.3300 0.4800 3.3900 0.5400 ;
        RECT 3.2250 0.1350 3.2850 0.1950 ;
        RECT 3.2250 0.8325 3.2850 0.8925 ;
        RECT 3.1200 0.4800 3.1800 0.5400 ;
        RECT 3.0150 0.3075 3.0750 0.3675 ;
        RECT 3.0150 0.6525 3.0750 0.7125 ;
        RECT 2.9100 0.4800 2.9700 0.5400 ;
        RECT 2.8050 0.1200 2.8650 0.1800 ;
        RECT 2.8050 0.8700 2.8650 0.9300 ;
        RECT 2.7000 0.4875 2.7600 0.5475 ;
        RECT 2.5950 0.7650 2.6550 0.8250 ;
        RECT 2.4900 0.4725 2.5500 0.5325 ;
        RECT 2.3850 0.2400 2.4450 0.3000 ;
        RECT 2.3850 0.8325 2.4450 0.8925 ;
        RECT 2.1750 0.2700 2.2350 0.3300 ;
        RECT 2.1750 0.7200 2.2350 0.7800 ;
        RECT 2.0700 0.4725 2.1300 0.5325 ;
        RECT 1.9650 0.1200 2.0250 0.1800 ;
        RECT 1.9650 0.8625 2.0250 0.9225 ;
        RECT 1.8675 0.4650 1.9275 0.5250 ;
        RECT 1.7550 0.2325 1.8150 0.2925 ;
        RECT 1.7550 0.6525 1.8150 0.7125 ;
        RECT 1.5450 0.1575 1.6050 0.2175 ;
        RECT 1.5450 0.8325 1.6050 0.8925 ;
        RECT 1.4325 0.6450 1.4925 0.7050 ;
        RECT 1.3350 0.1275 1.3950 0.1875 ;
        RECT 1.3350 0.8700 1.3950 0.9300 ;
        RECT 1.2300 0.3150 1.2900 0.3750 ;
        RECT 1.0200 0.3525 1.0800 0.4125 ;
        RECT 1.0200 0.6150 1.0800 0.6750 ;
        RECT 0.9150 0.1575 0.9750 0.2175 ;
        RECT 0.9150 0.8325 0.9750 0.8925 ;
        RECT 0.8175 0.3975 0.8775 0.4575 ;
        RECT 0.7050 0.1575 0.7650 0.2175 ;
        RECT 0.7050 0.8100 0.7650 0.8700 ;
        RECT 0.6075 0.5775 0.6675 0.6375 ;
        RECT 0.4950 0.2100 0.5550 0.2700 ;
        RECT 0.4950 0.8100 0.5550 0.8700 ;
        RECT 0.3900 0.4650 0.4500 0.5250 ;
        RECT 0.2850 0.1200 0.3450 0.1800 ;
        RECT 0.1725 0.4650 0.2325 0.5250 ;
        RECT 0.0750 0.2100 0.1350 0.2700 ;
        RECT 0.0750 0.8325 0.1350 0.8925 ;
        LAYER M1 ;
        RECT 2.9175 0.4725 3.6450 0.5475 ;
        RECT 2.9925 0.2775 3.5175 0.3975 ;
        RECT 2.9925 0.6225 3.5175 0.7425 ;
        RECT 2.8425 0.2550 2.9175 0.7950 ;
        RECT 2.4525 0.2550 2.8425 0.3300 ;
        RECT 2.6775 0.7200 2.8425 0.7950 ;
        RECT 2.6250 0.4050 2.7675 0.6450 ;
        RECT 2.5725 0.7200 2.6775 0.8550 ;
        RECT 2.3925 0.4425 2.5500 0.5625 ;
        RECT 2.3775 0.2100 2.4525 0.3300 ;
        RECT 2.2275 0.4125 2.3925 0.5625 ;
        RECT 1.9950 0.2625 2.2650 0.3375 ;
        RECT 1.9950 0.7125 2.2650 0.7875 ;
        RECT 2.0700 0.4425 2.2275 0.5625 ;
        RECT 1.9200 0.2625 1.9950 0.7875 ;
        RECT 1.8675 0.4350 1.9200 0.5550 ;
        RECT 1.7925 0.2025 1.8375 0.3225 ;
        RECT 1.7925 0.6300 1.8375 0.7350 ;
        RECT 1.7175 0.2025 1.7925 0.7350 ;
        RECT 1.5675 0.1500 1.6425 0.9000 ;
        RECT 1.5150 0.1500 1.5675 0.3600 ;
        RECT 1.5150 0.8250 1.5675 0.9000 ;
        RECT 1.2975 0.2850 1.5150 0.3600 ;
        RECT 1.2600 0.6150 1.4925 0.7350 ;
        RECT 1.2225 0.2850 1.2975 0.4050 ;
        RECT 1.1850 0.6150 1.2600 0.9000 ;
        RECT 0.8850 0.8100 1.1850 0.9000 ;
        RECT 1.0200 0.3225 1.1400 0.4875 ;
        RECT 0.9150 0.5625 1.0800 0.7050 ;
        RECT 0.8175 0.3675 1.0200 0.4875 ;
        RECT 0.7425 0.1500 1.0125 0.2250 ;
        RECT 0.6975 0.6150 0.9150 0.7050 ;
        RECT 0.4875 0.7800 0.7800 0.9000 ;
        RECT 0.6675 0.1500 0.7425 0.5025 ;
        RECT 0.5775 0.5775 0.6975 0.7050 ;
        RECT 0.5775 0.4125 0.6675 0.5025 ;
        RECT 0.4875 0.1800 0.5625 0.3300 ;
        RECT 0.1425 0.2550 0.4875 0.3300 ;
        RECT 0.3075 0.4050 0.4725 0.6000 ;
        RECT 0.2475 0.6750 0.3825 0.8175 ;
        RECT 0.2325 0.6750 0.2475 0.7500 ;
        RECT 0.1575 0.4350 0.2325 0.7500 ;
        RECT 0.0675 0.1800 0.1425 0.3300 ;
        LAYER VIA1 ;
        RECT 2.6775 0.5250 2.7525 0.6000 ;
        RECT 1.9200 0.5625 1.9950 0.6375 ;
        RECT 1.7175 0.3675 1.7925 0.4425 ;
        RECT 1.5675 0.7125 1.6425 0.7875 ;
        RECT 1.1850 0.7125 1.2600 0.7875 ;
        RECT 1.0650 0.3675 1.1400 0.4425 ;
        RECT 0.9600 0.5625 1.0350 0.6375 ;
        RECT 0.6225 0.4275 0.6975 0.5025 ;
        LAYER M2 ;
        RECT 2.6625 0.4800 2.7675 0.7875 ;
        RECT 1.5225 0.7125 2.6625 0.7875 ;
        RECT 0.9150 0.5625 2.0400 0.6375 ;
        RECT 1.0200 0.3675 1.8375 0.4425 ;
        RECT 0.7650 0.7125 1.3050 0.7875 ;
        RECT 0.6900 0.4275 0.7650 0.7875 ;
        RECT 0.5775 0.4275 0.6900 0.5025 ;
    END
END CKLNQ_0111


MACRO CKLNQ_1010
    CLASS CORE ;
    FOREIGN CKLNQ_1010 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.1500 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN TE
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.0900 0.7125 0.5700 0.7875 ;
        VIA 0.3150 0.7500 VIA12_square ;
        END
    END TE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 3.0375 0.2025 3.1125 0.8325 ;
        RECT 3.0075 0.2025 3.0375 0.3225 ;
        RECT 3.0075 0.6675 3.0375 0.8325 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.4275 0.2625 0.8925 0.3375 ;
        RECT 0.3525 0.2625 0.4275 0.5400 ;
        VIA 0.3900 0.4575 VIA12_square ;
        END
    END E
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 2.0250 0.4125 2.5500 0.4875 ;
        VIA 2.3100 0.4500 VIA12_square ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 2.8950 -0.0750 3.1500 0.0750 ;
        RECT 2.7750 -0.0750 2.8950 0.1800 ;
        RECT 2.0550 -0.0750 2.7750 0.0750 ;
        RECT 1.9350 -0.0750 2.0550 0.1875 ;
        RECT 1.4250 -0.0750 1.9350 0.0750 ;
        RECT 1.3050 -0.0750 1.4250 0.2100 ;
        RECT 0.3750 -0.0750 1.3050 0.0750 ;
        RECT 0.2550 -0.0750 0.3750 0.1800 ;
        RECT 0.0000 -0.0750 0.2550 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 2.8950 0.9750 3.1500 1.1250 ;
        RECT 2.7750 0.8700 2.8950 1.1250 ;
        RECT 2.4750 0.9750 2.7750 1.1250 ;
        RECT 2.3700 0.8025 2.4750 1.1250 ;
        RECT 2.0550 0.9750 2.3700 1.1250 ;
        RECT 1.9350 0.8625 2.0550 1.1250 ;
        RECT 1.4100 0.9750 1.9350 1.1250 ;
        RECT 1.3350 0.8400 1.4100 1.1250 ;
        RECT 0.1650 0.9750 1.3350 1.1250 ;
        RECT 0.0450 0.8250 0.1650 1.1250 ;
        RECT 0.0000 0.9750 0.0450 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 3.0150 0.2325 3.0750 0.2925 ;
        RECT 3.0150 0.7425 3.0750 0.8025 ;
        RECT 2.9025 0.4950 2.9625 0.5550 ;
        RECT 2.8050 0.1200 2.8650 0.1800 ;
        RECT 2.8050 0.8700 2.8650 0.9300 ;
        RECT 2.7000 0.4875 2.7600 0.5475 ;
        RECT 2.5950 0.8100 2.6550 0.8700 ;
        RECT 2.4900 0.4725 2.5500 0.5325 ;
        RECT 2.3850 0.2250 2.4450 0.2850 ;
        RECT 2.3850 0.8325 2.4450 0.8925 ;
        RECT 2.1750 0.2700 2.2350 0.3300 ;
        RECT 2.1750 0.7200 2.2350 0.7800 ;
        RECT 2.0700 0.4725 2.1300 0.5325 ;
        RECT 1.9650 0.1200 2.0250 0.1800 ;
        RECT 1.9650 0.8625 2.0250 0.9225 ;
        RECT 1.8675 0.4650 1.9275 0.5250 ;
        RECT 1.7550 0.2325 1.8150 0.2925 ;
        RECT 1.7550 0.6525 1.8150 0.7125 ;
        RECT 1.5450 0.1575 1.6050 0.2175 ;
        RECT 1.5450 0.8325 1.6050 0.8925 ;
        RECT 1.4325 0.6450 1.4925 0.7050 ;
        RECT 1.3350 0.1275 1.3950 0.1875 ;
        RECT 1.3350 0.8700 1.3950 0.9300 ;
        RECT 1.2300 0.3150 1.2900 0.3750 ;
        RECT 1.0200 0.3525 1.0800 0.4125 ;
        RECT 1.0200 0.6150 1.0800 0.6750 ;
        RECT 0.9150 0.1575 0.9750 0.2175 ;
        RECT 0.9150 0.8325 0.9750 0.8925 ;
        RECT 0.8175 0.3975 0.8775 0.4575 ;
        RECT 0.7050 0.1575 0.7650 0.2175 ;
        RECT 0.7050 0.8100 0.7650 0.8700 ;
        RECT 0.6075 0.5775 0.6675 0.6375 ;
        RECT 0.4950 0.2100 0.5550 0.2700 ;
        RECT 0.4950 0.8100 0.5550 0.8700 ;
        RECT 0.3900 0.4650 0.4500 0.5250 ;
        RECT 0.2850 0.1200 0.3450 0.1800 ;
        RECT 0.1725 0.4650 0.2325 0.5250 ;
        RECT 0.0750 0.2100 0.1350 0.2700 ;
        RECT 0.0750 0.8325 0.1350 0.8925 ;
        LAYER M1 ;
        RECT 2.9175 0.4650 2.9625 0.5850 ;
        RECT 2.8425 0.2550 2.9175 0.7950 ;
        RECT 2.4525 0.2550 2.8425 0.3300 ;
        RECT 2.6775 0.7200 2.8425 0.7950 ;
        RECT 2.6250 0.4050 2.7675 0.6450 ;
        RECT 2.5725 0.7200 2.6775 0.8925 ;
        RECT 2.3925 0.4425 2.5500 0.5625 ;
        RECT 2.3775 0.1800 2.4525 0.3300 ;
        RECT 2.2275 0.4125 2.3925 0.5625 ;
        RECT 1.9950 0.2625 2.2650 0.3375 ;
        RECT 1.9950 0.7125 2.2650 0.7875 ;
        RECT 2.0700 0.4425 2.2275 0.5625 ;
        RECT 1.9200 0.2625 1.9950 0.7875 ;
        RECT 1.8675 0.4350 1.9200 0.5550 ;
        RECT 1.7925 0.2025 1.8375 0.3225 ;
        RECT 1.7925 0.6300 1.8375 0.7350 ;
        RECT 1.7175 0.2025 1.7925 0.7350 ;
        RECT 1.5675 0.1500 1.6425 0.9000 ;
        RECT 1.5150 0.1500 1.5675 0.3600 ;
        RECT 1.5150 0.8250 1.5675 0.9000 ;
        RECT 1.2975 0.2850 1.5150 0.3600 ;
        RECT 1.2600 0.6150 1.4925 0.7350 ;
        RECT 1.2225 0.2850 1.2975 0.4050 ;
        RECT 1.1850 0.6150 1.2600 0.9000 ;
        RECT 0.8850 0.8100 1.1850 0.9000 ;
        RECT 1.0200 0.3225 1.1400 0.4875 ;
        RECT 0.9150 0.5625 1.0800 0.7050 ;
        RECT 0.8175 0.3675 1.0200 0.4875 ;
        RECT 0.7425 0.1500 1.0125 0.2250 ;
        RECT 0.6975 0.6150 0.9150 0.7050 ;
        RECT 0.4875 0.7800 0.7800 0.9000 ;
        RECT 0.6675 0.1500 0.7425 0.5025 ;
        RECT 0.5775 0.5775 0.6975 0.7050 ;
        RECT 0.5775 0.4125 0.6675 0.5025 ;
        RECT 0.4875 0.1800 0.5625 0.3300 ;
        RECT 0.1425 0.2550 0.4875 0.3300 ;
        RECT 0.3075 0.4050 0.4725 0.6000 ;
        RECT 0.2475 0.6750 0.3825 0.8175 ;
        RECT 0.2325 0.6750 0.2475 0.7500 ;
        RECT 0.1575 0.4350 0.2325 0.7500 ;
        RECT 0.0675 0.1800 0.1425 0.3300 ;
        LAYER VIA1 ;
        RECT 2.6775 0.5250 2.7525 0.6000 ;
        RECT 1.9200 0.5625 1.9950 0.6375 ;
        RECT 1.7175 0.3675 1.7925 0.4425 ;
        RECT 1.5675 0.7125 1.6425 0.7875 ;
        RECT 1.1850 0.7125 1.2600 0.7875 ;
        RECT 1.0650 0.3675 1.1400 0.4425 ;
        RECT 0.9600 0.5625 1.0350 0.6375 ;
        RECT 0.6225 0.4275 0.6975 0.5025 ;
        LAYER M2 ;
        RECT 2.6775 0.4800 2.7525 0.7875 ;
        RECT 1.5225 0.7125 2.6775 0.7875 ;
        RECT 0.9150 0.5625 2.0400 0.6375 ;
        RECT 1.0200 0.3675 1.8375 0.4425 ;
        RECT 0.7650 0.7125 1.3050 0.7875 ;
        RECT 0.6900 0.4275 0.7650 0.7875 ;
        RECT 0.5775 0.4275 0.6900 0.5025 ;
    END
END CKLNQ_1010


MACRO CKLNQ_1100
    CLASS CORE ;
    FOREIGN CKLNQ_1100 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.5600 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN TE
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.0900 0.7125 0.5700 0.7875 ;
        VIA 0.3150 0.7500 VIA12_square ;
        END
    END TE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 5.9325 0.2775 6.0900 0.3975 ;
        RECT 5.9325 0.6225 6.0900 0.7425 ;
        RECT 5.6175 0.2775 5.9325 0.7425 ;
        RECT 5.4600 0.2775 5.6175 0.3975 ;
        RECT 5.4600 0.6225 5.6175 0.7425 ;
        VIA 5.9325 0.3375 VIA12_slot ;
        VIA 5.9325 0.6825 VIA12_slot ;
        VIA 5.6175 0.3375 VIA12_slot ;
        VIA 5.6175 0.6825 VIA12_slot ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.4275 0.2625 0.8925 0.3375 ;
        RECT 0.3525 0.2625 0.4275 0.5400 ;
        VIA 0.3900 0.4575 VIA12_square ;
        END
    END E
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 3.6375 0.2625 3.7125 0.5925 ;
        RECT 2.8650 0.2625 3.6375 0.3375 ;
        RECT 2.8650 0.4650 2.9700 0.5400 ;
        RECT 2.7900 0.1650 2.8650 0.5400 ;
        RECT 2.2650 0.1650 2.7900 0.2400 ;
        RECT 2.1900 0.1650 2.2650 0.4800 ;
        RECT 2.0700 0.4050 2.1900 0.4800 ;
        VIA 3.6750 0.5100 VIA12_square ;
        VIA 2.8725 0.5025 VIA12_square ;
        VIA 2.1525 0.4425 VIA12_square ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 7.4925 -0.0750 7.5600 0.0750 ;
        RECT 7.4175 -0.0750 7.4925 0.2925 ;
        RECT 7.0950 -0.0750 7.4175 0.0750 ;
        RECT 6.9750 -0.0750 7.0950 0.2025 ;
        RECT 6.6750 -0.0750 6.9750 0.0750 ;
        RECT 6.5550 -0.0750 6.6750 0.2025 ;
        RECT 6.2550 -0.0750 6.5550 0.0750 ;
        RECT 6.1350 -0.0750 6.2550 0.2025 ;
        RECT 5.8350 -0.0750 6.1350 0.0750 ;
        RECT 5.7150 -0.0750 5.8350 0.2025 ;
        RECT 5.4150 -0.0750 5.7150 0.0750 ;
        RECT 5.2950 -0.0750 5.4150 0.2025 ;
        RECT 4.9950 -0.0750 5.2950 0.0750 ;
        RECT 4.8750 -0.0750 4.9950 0.2025 ;
        RECT 4.5750 -0.0750 4.8750 0.0750 ;
        RECT 4.4550 -0.0750 4.5750 0.2025 ;
        RECT 4.1550 -0.0750 4.4550 0.0750 ;
        RECT 4.0500 -0.0750 4.1550 0.2250 ;
        RECT 3.3150 -0.0750 4.0500 0.0750 ;
        RECT 3.1950 -0.0750 3.3150 0.2025 ;
        RECT 2.4600 -0.0750 3.1950 0.0750 ;
        RECT 2.3550 -0.0750 2.4600 0.2475 ;
        RECT 2.0550 -0.0750 2.3550 0.0750 ;
        RECT 1.9350 -0.0750 2.0550 0.1800 ;
        RECT 1.4250 -0.0750 1.9350 0.0750 ;
        RECT 1.3050 -0.0750 1.4250 0.2100 ;
        RECT 0.3750 -0.0750 1.3050 0.0750 ;
        RECT 0.2550 -0.0750 0.3750 0.1800 ;
        RECT 0.0000 -0.0750 0.2550 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 7.5075 0.9750 7.5600 1.1250 ;
        RECT 7.4025 0.6450 7.5075 1.1250 ;
        RECT 7.0950 0.9750 7.4025 1.1250 ;
        RECT 6.9750 0.8250 7.0950 1.1250 ;
        RECT 6.6750 0.9750 6.9750 1.1250 ;
        RECT 6.5550 0.8250 6.6750 1.1250 ;
        RECT 6.2550 0.9750 6.5550 1.1250 ;
        RECT 6.1350 0.8250 6.2550 1.1250 ;
        RECT 5.8350 0.9750 6.1350 1.1250 ;
        RECT 5.7150 0.8250 5.8350 1.1250 ;
        RECT 5.4150 0.9750 5.7150 1.1250 ;
        RECT 5.2950 0.8250 5.4150 1.1250 ;
        RECT 4.9950 0.9750 5.2950 1.1250 ;
        RECT 4.8750 0.8250 4.9950 1.1250 ;
        RECT 4.5750 0.9750 4.8750 1.1250 ;
        RECT 4.4550 0.8250 4.5750 1.1250 ;
        RECT 4.1550 0.9750 4.4550 1.1250 ;
        RECT 4.0350 0.8700 4.1550 1.1250 ;
        RECT 3.7350 0.9750 4.0350 1.1250 ;
        RECT 3.6150 0.8700 3.7350 1.1250 ;
        RECT 3.3150 0.9750 3.6150 1.1250 ;
        RECT 3.1950 0.8475 3.3150 1.1250 ;
        RECT 2.8950 0.9750 3.1950 1.1250 ;
        RECT 2.7750 0.8475 2.8950 1.1250 ;
        RECT 2.4525 0.9750 2.7750 1.1250 ;
        RECT 2.3775 0.8025 2.4525 1.1250 ;
        RECT 2.0550 0.9750 2.3775 1.1250 ;
        RECT 1.9350 0.8625 2.0550 1.1250 ;
        RECT 1.4100 0.9750 1.9350 1.1250 ;
        RECT 1.3350 0.8400 1.4100 1.1250 ;
        RECT 0.1650 0.9750 1.3350 1.1250 ;
        RECT 0.0450 0.8250 0.1650 1.1250 ;
        RECT 0.0000 0.9750 0.0450 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 7.4250 0.2025 7.4850 0.2625 ;
        RECT 7.4250 0.6675 7.4850 0.7275 ;
        RECT 7.4250 0.8325 7.4850 0.8925 ;
        RECT 7.3200 0.4800 7.3800 0.5400 ;
        RECT 7.2150 0.3075 7.2750 0.3675 ;
        RECT 7.2150 0.6525 7.2750 0.7125 ;
        RECT 7.1100 0.4800 7.1700 0.5400 ;
        RECT 7.0050 0.1350 7.0650 0.1950 ;
        RECT 7.0050 0.8325 7.0650 0.8925 ;
        RECT 6.9000 0.4800 6.9600 0.5400 ;
        RECT 6.7950 0.3075 6.8550 0.3675 ;
        RECT 6.7950 0.6525 6.8550 0.7125 ;
        RECT 6.6900 0.4800 6.7500 0.5400 ;
        RECT 6.5850 0.1350 6.6450 0.1950 ;
        RECT 6.5850 0.8325 6.6450 0.8925 ;
        RECT 6.4800 0.4800 6.5400 0.5400 ;
        RECT 6.3750 0.3075 6.4350 0.3675 ;
        RECT 6.3750 0.6525 6.4350 0.7125 ;
        RECT 6.2700 0.4800 6.3300 0.5400 ;
        RECT 6.1650 0.1350 6.2250 0.1950 ;
        RECT 6.1650 0.8325 6.2250 0.8925 ;
        RECT 6.0600 0.4800 6.1200 0.5400 ;
        RECT 5.9550 0.3075 6.0150 0.3675 ;
        RECT 5.9550 0.6525 6.0150 0.7125 ;
        RECT 5.8500 0.4800 5.9100 0.5400 ;
        RECT 5.7450 0.1350 5.8050 0.1950 ;
        RECT 5.7450 0.8325 5.8050 0.8925 ;
        RECT 5.6400 0.4800 5.7000 0.5400 ;
        RECT 5.5350 0.3075 5.5950 0.3675 ;
        RECT 5.5350 0.6525 5.5950 0.7125 ;
        RECT 5.4300 0.4800 5.4900 0.5400 ;
        RECT 5.3250 0.1350 5.3850 0.1950 ;
        RECT 5.3250 0.8325 5.3850 0.8925 ;
        RECT 5.2200 0.4800 5.2800 0.5400 ;
        RECT 5.1150 0.3075 5.1750 0.3675 ;
        RECT 5.1150 0.6525 5.1750 0.7125 ;
        RECT 5.0100 0.4800 5.0700 0.5400 ;
        RECT 4.9050 0.1350 4.9650 0.1950 ;
        RECT 4.9050 0.8325 4.9650 0.8925 ;
        RECT 4.8000 0.4800 4.8600 0.5400 ;
        RECT 4.6950 0.3075 4.7550 0.3675 ;
        RECT 4.6950 0.6525 4.7550 0.7125 ;
        RECT 4.5900 0.4800 4.6500 0.5400 ;
        RECT 4.4850 0.1350 4.5450 0.1950 ;
        RECT 4.4850 0.8325 4.5450 0.8925 ;
        RECT 4.3800 0.4800 4.4400 0.5400 ;
        RECT 4.2750 0.3075 4.3350 0.3675 ;
        RECT 4.2750 0.6525 4.3350 0.7125 ;
        RECT 4.1700 0.4800 4.2300 0.5400 ;
        RECT 4.0650 0.1350 4.1250 0.1950 ;
        RECT 4.0650 0.8700 4.1250 0.9300 ;
        RECT 3.9600 0.4950 4.0200 0.5550 ;
        RECT 3.8550 0.1575 3.9150 0.2175 ;
        RECT 3.8550 0.7950 3.9150 0.8550 ;
        RECT 3.7500 0.4875 3.8100 0.5475 ;
        RECT 3.6450 0.3075 3.7050 0.3675 ;
        RECT 3.6450 0.8700 3.7050 0.9300 ;
        RECT 3.5400 0.4875 3.6000 0.5475 ;
        RECT 3.4350 0.2250 3.4950 0.2850 ;
        RECT 3.4350 0.8025 3.4950 0.8625 ;
        RECT 3.3300 0.4875 3.3900 0.5475 ;
        RECT 3.2250 0.1350 3.2850 0.1950 ;
        RECT 3.2250 0.8550 3.2850 0.9150 ;
        RECT 3.1200 0.4875 3.1800 0.5475 ;
        RECT 3.0150 0.2250 3.0750 0.2850 ;
        RECT 3.0150 0.8025 3.0750 0.8625 ;
        RECT 2.9100 0.4875 2.9700 0.5475 ;
        RECT 2.8050 0.3075 2.8650 0.3675 ;
        RECT 2.8050 0.8550 2.8650 0.9150 ;
        RECT 2.7000 0.4875 2.7600 0.5475 ;
        RECT 2.5950 0.1575 2.6550 0.2175 ;
        RECT 2.5950 0.8025 2.6550 0.8625 ;
        RECT 2.4900 0.4875 2.5500 0.5475 ;
        RECT 2.3850 0.1575 2.4450 0.2175 ;
        RECT 2.3850 0.8325 2.4450 0.8925 ;
        RECT 2.1750 0.2175 2.2350 0.2775 ;
        RECT 2.1750 0.7650 2.2350 0.8250 ;
        RECT 2.0700 0.4725 2.1300 0.5325 ;
        RECT 1.9650 0.1200 2.0250 0.1800 ;
        RECT 1.9650 0.8625 2.0250 0.9225 ;
        RECT 1.8675 0.4650 1.9275 0.5250 ;
        RECT 1.7550 0.2325 1.8150 0.2925 ;
        RECT 1.7550 0.6525 1.8150 0.7125 ;
        RECT 1.5450 0.1575 1.6050 0.2175 ;
        RECT 1.5450 0.8325 1.6050 0.8925 ;
        RECT 1.4325 0.6450 1.4925 0.7050 ;
        RECT 1.3350 0.1275 1.3950 0.1875 ;
        RECT 1.3350 0.8700 1.3950 0.9300 ;
        RECT 1.2300 0.3150 1.2900 0.3750 ;
        RECT 1.0200 0.3525 1.0800 0.4125 ;
        RECT 1.0200 0.6150 1.0800 0.6750 ;
        RECT 0.9150 0.1575 0.9750 0.2175 ;
        RECT 0.9150 0.8325 0.9750 0.8925 ;
        RECT 0.8175 0.3975 0.8775 0.4575 ;
        RECT 0.7050 0.1575 0.7650 0.2175 ;
        RECT 0.7050 0.8100 0.7650 0.8700 ;
        RECT 0.6075 0.5775 0.6675 0.6375 ;
        RECT 0.4950 0.2100 0.5550 0.2700 ;
        RECT 0.4950 0.8100 0.5550 0.8700 ;
        RECT 0.3900 0.4650 0.4500 0.5250 ;
        RECT 0.2850 0.1200 0.3450 0.1800 ;
        RECT 0.1725 0.4650 0.2325 0.5250 ;
        RECT 0.0750 0.2100 0.1350 0.2700 ;
        RECT 0.0750 0.8325 0.1350 0.8925 ;
        LAYER M1 ;
        RECT 4.2000 0.4725 7.4100 0.5475 ;
        RECT 4.2750 0.2775 7.3050 0.3975 ;
        RECT 4.2750 0.6225 7.3050 0.7425 ;
        RECT 4.1250 0.3000 4.2000 0.7950 ;
        RECT 3.6150 0.3000 4.1250 0.3750 ;
        RECT 3.9450 0.7200 4.1250 0.7950 ;
        RECT 3.8850 0.4500 4.0500 0.6450 ;
        RECT 3.5025 0.1500 3.9450 0.2250 ;
        RECT 3.8250 0.7200 3.9450 0.8700 ;
        RECT 3.5250 0.7200 3.8250 0.7950 ;
        RECT 3.5325 0.4500 3.8100 0.5775 ;
        RECT 3.4050 0.6975 3.5250 0.8775 ;
        RECT 3.4275 0.1500 3.5025 0.3525 ;
        RECT 3.0825 0.2775 3.4275 0.3525 ;
        RECT 3.1050 0.6975 3.4050 0.7725 ;
        RECT 3.1200 0.4500 3.3900 0.5775 ;
        RECT 2.9850 0.6975 3.1050 0.8775 ;
        RECT 3.0075 0.1500 3.0825 0.3525 ;
        RECT 2.5650 0.1500 3.0075 0.2250 ;
        RECT 2.8725 0.6975 2.9850 0.7725 ;
        RECT 2.7000 0.4500 2.9700 0.5775 ;
        RECT 2.6250 0.3000 2.8950 0.3750 ;
        RECT 2.7000 0.6525 2.8725 0.7725 ;
        RECT 2.6850 0.6975 2.7000 0.7725 ;
        RECT 2.5650 0.6975 2.6850 0.8775 ;
        RECT 2.5650 0.3000 2.6250 0.3975 ;
        RECT 2.3775 0.4725 2.6250 0.6075 ;
        RECT 2.4300 0.3225 2.5650 0.3975 ;
        RECT 2.1600 0.1875 2.2350 0.3300 ;
        RECT 2.0700 0.4050 2.2350 0.6000 ;
        RECT 2.1600 0.7125 2.2350 0.8550 ;
        RECT 1.9950 0.2550 2.1600 0.3300 ;
        RECT 1.9950 0.7125 2.1600 0.7875 ;
        RECT 1.9200 0.2550 1.9950 0.7875 ;
        RECT 1.8675 0.4350 1.9200 0.5550 ;
        RECT 1.7925 0.2025 1.8375 0.3225 ;
        RECT 1.7925 0.6300 1.8375 0.7350 ;
        RECT 1.7175 0.2025 1.7925 0.7350 ;
        RECT 1.5675 0.1500 1.6425 0.9000 ;
        RECT 1.5150 0.1500 1.5675 0.3600 ;
        RECT 1.5150 0.8250 1.5675 0.9000 ;
        RECT 1.2975 0.2850 1.5150 0.3600 ;
        RECT 1.2600 0.6150 1.4925 0.7350 ;
        RECT 1.2225 0.2850 1.2975 0.4050 ;
        RECT 1.1850 0.6150 1.2600 0.9000 ;
        RECT 0.8850 0.8100 1.1850 0.9000 ;
        RECT 1.0200 0.3225 1.1400 0.4875 ;
        RECT 0.9150 0.5625 1.0800 0.7050 ;
        RECT 0.8175 0.3675 1.0200 0.4875 ;
        RECT 0.7425 0.1500 1.0125 0.2250 ;
        RECT 0.6975 0.6150 0.9150 0.7050 ;
        RECT 0.4875 0.7800 0.7800 0.9000 ;
        RECT 0.6675 0.1500 0.7425 0.5025 ;
        RECT 0.5775 0.5775 0.6975 0.7050 ;
        RECT 0.5775 0.4125 0.6675 0.5025 ;
        RECT 0.4875 0.1800 0.5625 0.3300 ;
        RECT 0.1425 0.2550 0.4875 0.3300 ;
        RECT 0.3075 0.4050 0.4725 0.6000 ;
        RECT 0.2475 0.6750 0.3825 0.8175 ;
        RECT 0.2325 0.6750 0.2475 0.7500 ;
        RECT 0.1575 0.4350 0.2325 0.7500 ;
        RECT 0.0675 0.1800 0.1425 0.3300 ;
        LAYER VIA1 ;
        RECT 3.9375 0.4950 4.0125 0.5700 ;
        RECT 3.2250 0.5025 3.3000 0.5775 ;
        RECT 2.7525 0.6600 2.8275 0.7350 ;
        RECT 2.4900 0.3225 2.5650 0.3975 ;
        RECT 2.4300 0.5175 2.5050 0.5925 ;
        RECT 1.9200 0.5625 1.9950 0.6375 ;
        RECT 1.7175 0.3675 1.7925 0.4425 ;
        RECT 1.5675 0.7125 1.6425 0.7875 ;
        RECT 1.1850 0.7125 1.2600 0.7875 ;
        RECT 1.0650 0.3675 1.1400 0.4425 ;
        RECT 0.9600 0.5625 1.0350 0.6375 ;
        RECT 0.6225 0.4275 0.6975 0.5025 ;
        LAYER M2 ;
        RECT 5.9625 0.2775 6.0900 0.3975 ;
        RECT 5.9625 0.6225 6.0900 0.7425 ;
        RECT 5.4600 0.2775 5.5875 0.3975 ;
        RECT 5.4600 0.6225 5.5875 0.7425 ;
        RECT 3.9375 0.4500 4.0125 0.8850 ;
        RECT 3.3150 0.8100 3.9375 0.8850 ;
        RECT 3.2100 0.4575 3.3150 0.8850 ;
        RECT 2.5500 0.8100 3.2100 0.8850 ;
        RECT 2.7000 0.6600 2.8725 0.7350 ;
        RECT 2.6250 0.3225 2.7000 0.7350 ;
        RECT 2.4450 0.3225 2.6250 0.3975 ;
        RECT 2.4750 0.5025 2.5500 0.8850 ;
        RECT 2.3850 0.5025 2.4750 0.6075 ;
        RECT 1.5225 0.7125 2.4750 0.7875 ;
        RECT 0.9150 0.5625 2.0400 0.6375 ;
        RECT 1.0200 0.3675 1.8375 0.4425 ;
        RECT 0.7650 0.7125 1.3050 0.7875 ;
        RECT 0.6900 0.4275 0.7650 0.7875 ;
        RECT 0.5775 0.4275 0.6900 0.5025 ;
    END
END CKLNQ_1100


MACRO CKMUX2_0011
    CLASS CORE ;
    FOREIGN CKMUX2_0011 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.6800 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 1.5675 0.3000 1.6425 0.7425 ;
        RECT 1.4025 0.3000 1.5675 0.3750 ;
        RECT 1.4025 0.6675 1.5675 0.7425 ;
        RECT 1.3275 0.2025 1.4025 0.3750 ;
        RECT 1.3275 0.6675 1.4025 0.8325 ;
        END
    END Z
    PIN S
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.5025 0.7125 0.9225 0.7875 ;
        RECT 0.3975 0.4875 0.5025 0.7875 ;
        VIA 0.4500 0.5625 VIA12_square ;
        END
    END S
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.6525 0.4125 1.1175 0.4875 ;
        VIA 1.0200 0.4500 VIA12_square ;
        END
    END I1
    PIN I0
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.4275 0.2625 0.8925 0.3375 ;
        VIA 0.5625 0.3000 VIA12_square ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.6350 -0.0750 1.6800 0.0750 ;
        RECT 1.5150 -0.0750 1.6350 0.2250 ;
        RECT 1.2150 -0.0750 1.5150 0.0750 ;
        RECT 1.0950 -0.0750 1.2150 0.1800 ;
        RECT 0.3750 -0.0750 1.0950 0.0750 ;
        RECT 0.2550 -0.0750 0.3750 0.1800 ;
        RECT 0.0000 -0.0750 0.2550 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.6350 0.9750 1.6800 1.1250 ;
        RECT 1.5150 0.8250 1.6350 1.1250 ;
        RECT 1.2300 0.9750 1.5150 1.1250 ;
        RECT 1.1250 0.8400 1.2300 1.1250 ;
        RECT 0.3750 0.9750 1.1250 1.1250 ;
        RECT 0.2550 0.8625 0.3750 1.1250 ;
        RECT 0.0000 0.9750 0.2550 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.5450 0.1575 1.6050 0.2175 ;
        RECT 1.5450 0.8325 1.6050 0.8925 ;
        RECT 1.4325 0.4800 1.4925 0.5400 ;
        RECT 1.3350 0.2325 1.3950 0.2925 ;
        RECT 1.3350 0.7200 1.3950 0.7800 ;
        RECT 1.2300 0.4800 1.2900 0.5400 ;
        RECT 1.1250 0.1200 1.1850 0.1800 ;
        RECT 1.1250 0.8700 1.1850 0.9300 ;
        RECT 1.0200 0.4875 1.0800 0.5475 ;
        RECT 0.8100 0.6375 0.8700 0.6975 ;
        RECT 0.8025 0.3900 0.8625 0.4500 ;
        RECT 0.7050 0.1725 0.7650 0.2325 ;
        RECT 0.7050 0.8325 0.7650 0.8925 ;
        RECT 0.5925 0.3450 0.6525 0.4050 ;
        RECT 0.3825 0.3150 0.4425 0.3750 ;
        RECT 0.3825 0.5550 0.4425 0.6150 ;
        RECT 0.2850 0.1200 0.3450 0.1800 ;
        RECT 0.2850 0.8700 0.3450 0.9300 ;
        RECT 0.0750 0.7950 0.1350 0.8550 ;
        RECT 0.1875 0.5250 0.2475 0.5850 ;
        RECT 0.0750 0.1575 0.1350 0.2175 ;
        LAYER M1 ;
        RECT 1.2525 0.4500 1.4925 0.5700 ;
        RECT 1.1775 0.2550 1.2525 0.7650 ;
        RECT 1.0200 0.2550 1.1775 0.3300 ;
        RECT 1.0500 0.6900 1.1775 0.7650 ;
        RECT 0.9750 0.4050 1.1025 0.6150 ;
        RECT 0.9750 0.6900 1.0500 0.9000 ;
        RECT 0.9450 0.1500 1.0200 0.3300 ;
        RECT 0.9375 0.4050 0.9750 0.5400 ;
        RECT 0.6750 0.8250 0.9750 0.9000 ;
        RECT 0.6825 0.1500 0.9450 0.2550 ;
        RECT 0.7800 0.6375 0.9000 0.7500 ;
        RECT 0.7875 0.3600 0.8625 0.5625 ;
        RECT 0.6525 0.4875 0.7875 0.5625 ;
        RECT 0.6150 0.6750 0.7800 0.7500 ;
        RECT 0.6075 0.3300 0.6825 0.4125 ;
        RECT 0.5850 0.4875 0.6525 0.6000 ;
        RECT 0.5475 0.6750 0.6150 0.7650 ;
        RECT 0.5175 0.1500 0.6075 0.4125 ;
        RECT 0.4725 0.5250 0.5850 0.6000 ;
        RECT 0.1425 0.6900 0.5475 0.7650 ;
        RECT 0.4875 0.1500 0.5175 0.2250 ;
        RECT 0.2925 0.5250 0.4725 0.6150 ;
        RECT 0.3375 0.2850 0.4425 0.4050 ;
        RECT 0.1650 0.3300 0.3375 0.4050 ;
        RECT 0.1875 0.4800 0.2925 0.6150 ;
        RECT 0.1125 0.1500 0.1650 0.4050 ;
        RECT 0.1125 0.6900 0.1425 0.9000 ;
        RECT 0.0375 0.1500 0.1125 0.9000 ;
    END
END CKMUX2_0011


MACRO CKMUX2_0111
    CLASS CORE ;
    FOREIGN CKMUX2_0111 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.7300 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 2.0475 0.2625 2.3625 0.7725 ;
        VIA 2.2050 0.3225 VIA12_slot ;
        VIA 2.2050 0.7125 VIA12_slot ;
        END
    END Z
    PIN S
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.8550 0.3375 0.9900 0.4875 ;
        RECT 0.6750 0.4125 0.8550 0.4875 ;
        RECT 0.6000 0.4125 0.6750 0.6375 ;
        RECT 0.1200 0.5625 0.6000 0.6375 ;
        VIA 0.9225 0.4050 VIA12_square ;
        VIA 0.3675 0.6000 VIA12_square ;
        END
    END S
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.6650 0.8625 1.9800 0.9375 ;
        RECT 1.5900 0.4125 1.6650 0.9375 ;
        RECT 1.2750 0.4125 1.5900 0.4875 ;
        VIA 1.6275 0.5025 VIA12_square ;
        END
    END I1
    PIN I0
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.5700 0.1125 0.7275 0.1875 ;
        RECT 0.4650 0.1125 0.5700 0.2850 ;
        RECT 0.1125 0.1125 0.4650 0.1875 ;
        VIA 0.5175 0.2025 VIA12_square ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 2.6625 -0.0750 2.7300 0.0750 ;
        RECT 2.5875 -0.0750 2.6625 0.2625 ;
        RECT 2.2650 -0.0750 2.5875 0.0750 ;
        RECT 2.1450 -0.0750 2.2650 0.1950 ;
        RECT 1.8225 -0.0750 2.1450 0.0750 ;
        RECT 1.7475 -0.0750 1.8225 0.2475 ;
        RECT 1.4250 -0.0750 1.7475 0.0750 ;
        RECT 1.3050 -0.0750 1.4250 0.2250 ;
        RECT 0.3525 -0.0750 1.3050 0.0750 ;
        RECT 0.2775 -0.0750 0.3525 0.2100 ;
        RECT 0.0000 -0.0750 0.2775 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 2.6775 0.9750 2.7300 1.1250 ;
        RECT 2.5725 0.6375 2.6775 1.1250 ;
        RECT 2.2650 0.9750 2.5725 1.1250 ;
        RECT 2.1450 0.8400 2.2650 1.1250 ;
        RECT 1.8450 0.9750 2.1450 1.1250 ;
        RECT 1.7250 0.6975 1.8450 1.1250 ;
        RECT 1.4175 0.9750 1.7250 1.1250 ;
        RECT 1.3125 0.7800 1.4175 1.1250 ;
        RECT 0.3600 0.9750 1.3125 1.1250 ;
        RECT 0.2850 0.7950 0.3600 1.1250 ;
        RECT 0.0000 0.9750 0.2850 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 2.5950 0.1725 2.6550 0.2325 ;
        RECT 2.5950 0.6675 2.6550 0.7275 ;
        RECT 2.5950 0.8325 2.6550 0.8925 ;
        RECT 2.4900 0.4800 2.5500 0.5400 ;
        RECT 2.3850 0.2925 2.4450 0.3525 ;
        RECT 2.3850 0.6825 2.4450 0.7425 ;
        RECT 2.2800 0.4800 2.3400 0.5400 ;
        RECT 2.1750 0.1275 2.2350 0.1875 ;
        RECT 2.1750 0.8550 2.2350 0.9150 ;
        RECT 2.0700 0.4800 2.1300 0.5400 ;
        RECT 1.9650 0.2925 2.0250 0.3525 ;
        RECT 1.9650 0.6825 2.0250 0.7425 ;
        RECT 1.8600 0.4800 1.9200 0.5400 ;
        RECT 1.7550 0.1575 1.8150 0.2175 ;
        RECT 1.7550 0.7050 1.8150 0.7650 ;
        RECT 1.7550 0.8700 1.8150 0.9300 ;
        RECT 1.6425 0.4725 1.7025 0.5325 ;
        RECT 1.5450 0.1800 1.6050 0.2400 ;
        RECT 1.5450 0.7275 1.6050 0.7875 ;
        RECT 1.4400 0.4725 1.5000 0.5325 ;
        RECT 1.3350 0.1575 1.3950 0.2175 ;
        RECT 1.3350 0.8025 1.3950 0.8625 ;
        RECT 1.1250 0.1800 1.1850 0.2400 ;
        RECT 1.1250 0.8100 1.1850 0.8700 ;
        RECT 1.0200 0.3600 1.0800 0.4200 ;
        RECT 1.0200 0.6000 1.0800 0.6600 ;
        RECT 0.9150 0.1650 0.9750 0.2250 ;
        RECT 0.9150 0.8175 0.9750 0.8775 ;
        RECT 0.7050 0.1725 0.7650 0.2325 ;
        RECT 0.7050 0.8175 0.7650 0.8775 ;
        RECT 0.6000 0.4950 0.6600 0.5550 ;
        RECT 0.3900 0.3600 0.4500 0.4200 ;
        RECT 0.3900 0.6000 0.4500 0.6600 ;
        RECT 0.2850 0.1200 0.3450 0.1800 ;
        RECT 0.2850 0.8250 0.3450 0.8850 ;
        RECT 0.1875 0.5550 0.2475 0.6150 ;
        RECT 0.0750 0.1575 0.1350 0.2175 ;
        RECT 0.0750 0.7725 0.1350 0.8325 ;
        LAYER M1 ;
        RECT 1.8000 0.4575 2.5875 0.5625 ;
        RECT 1.9350 0.2700 2.4750 0.3750 ;
        RECT 1.9350 0.6600 2.4675 0.7650 ;
        RECT 1.4175 0.4500 1.7250 0.5550 ;
        RECT 1.5150 0.1725 1.6350 0.3750 ;
        RECT 1.5375 0.6300 1.6125 0.8175 ;
        RECT 1.2375 0.6300 1.5375 0.7050 ;
        RECT 1.2300 0.3000 1.5150 0.3750 ;
        RECT 1.1625 0.6300 1.2375 0.9000 ;
        RECT 1.1550 0.1500 1.2300 0.3750 ;
        RECT 1.1250 0.7800 1.1625 0.9000 ;
        RECT 1.1250 0.1500 1.1550 0.2700 ;
        RECT 0.8700 0.5550 1.0875 0.7050 ;
        RECT 0.8700 0.3300 1.0800 0.4800 ;
        RECT 0.6825 0.1500 1.0500 0.2550 ;
        RECT 0.6825 0.7950 1.0500 0.9000 ;
        RECT 0.6075 0.4875 0.7050 0.5625 ;
        RECT 0.5250 0.1500 0.6075 0.5625 ;
        RECT 0.4275 0.1500 0.5250 0.2550 ;
        RECT 0.3150 0.3300 0.4500 0.4500 ;
        RECT 0.3450 0.5250 0.4500 0.6900 ;
        RECT 0.1875 0.5250 0.3450 0.6450 ;
        RECT 0.1650 0.3300 0.3150 0.4050 ;
        RECT 0.1125 0.7275 0.2100 0.9000 ;
        RECT 0.1125 0.1500 0.1650 0.4050 ;
        RECT 0.0375 0.1500 0.1125 0.9000 ;
        LAYER VIA1 ;
        RECT 1.8375 0.4725 1.9125 0.5475 ;
        RECT 0.9375 0.1650 1.0125 0.2400 ;
        RECT 0.9375 0.8100 1.0125 0.8850 ;
        RECT 0.8850 0.5925 0.9600 0.6675 ;
        RECT 0.1350 0.7725 0.2100 0.8475 ;
        LAYER M2 ;
        RECT 1.8825 0.4275 1.9275 0.5925 ;
        RECT 1.8075 0.2625 1.8825 0.5925 ;
        RECT 1.1550 0.2625 1.8075 0.3375 ;
        RECT 1.0800 0.1500 1.1550 0.8700 ;
        RECT 0.9000 0.1500 1.0800 0.2550 ;
        RECT 1.0500 0.7950 1.0800 0.8700 ;
        RECT 0.9000 0.7950 1.0500 0.9000 ;
        RECT 0.8250 0.5775 0.9975 0.6825 ;
        RECT 0.7500 0.5775 0.8250 0.8475 ;
        RECT 0.0900 0.7725 0.7500 0.8475 ;
    END
END CKMUX2_0111


MACRO CKMUX2_1000
    CLASS CORE ;
    FOREIGN CKMUX2_1000 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.4700 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 1.3575 0.1500 1.4325 0.9000 ;
        RECT 1.3275 0.1500 1.3575 0.3825 ;
        RECT 1.3275 0.6675 1.3575 0.9000 ;
        END
    END Z
    PIN S
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.5025 0.7125 0.9225 0.7875 ;
        RECT 0.3975 0.4875 0.5025 0.7875 ;
        VIA 0.4500 0.5625 VIA12_square ;
        END
    END S
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.6525 0.4125 1.1175 0.4875 ;
        VIA 1.0200 0.4500 VIA12_square ;
        END
    END I1
    PIN I0
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.4275 0.2625 0.8925 0.3375 ;
        VIA 0.5625 0.3000 VIA12_square ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.2150 -0.0750 1.4700 0.0750 ;
        RECT 1.0950 -0.0750 1.2150 0.1800 ;
        RECT 0.3750 -0.0750 1.0950 0.0750 ;
        RECT 0.2550 -0.0750 0.3750 0.2100 ;
        RECT 0.0000 -0.0750 0.2550 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.2300 0.9750 1.4700 1.1250 ;
        RECT 1.1250 0.8400 1.2300 1.1250 ;
        RECT 0.3750 0.9750 1.1250 1.1250 ;
        RECT 0.2550 0.8400 0.3750 1.1250 ;
        RECT 0.0000 0.9750 0.2550 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.3350 0.1800 1.3950 0.2400 ;
        RECT 1.3350 0.8100 1.3950 0.8700 ;
        RECT 1.2225 0.4800 1.2825 0.5400 ;
        RECT 1.1250 0.1200 1.1850 0.1800 ;
        RECT 1.1250 0.8700 1.1850 0.9300 ;
        RECT 1.0200 0.4875 1.0800 0.5475 ;
        RECT 0.8100 0.6375 0.8700 0.6975 ;
        RECT 0.8025 0.3900 0.8625 0.4500 ;
        RECT 0.7050 0.1725 0.7650 0.2325 ;
        RECT 0.7050 0.8325 0.7650 0.8925 ;
        RECT 0.5925 0.3450 0.6525 0.4050 ;
        RECT 0.3825 0.3150 0.4425 0.3750 ;
        RECT 0.2850 0.8475 0.3450 0.9075 ;
        RECT 0.1875 0.5250 0.2475 0.5850 ;
        RECT 0.0750 0.1575 0.1350 0.2175 ;
        RECT 0.0750 0.8175 0.1350 0.8775 ;
        RECT 0.3825 0.5550 0.4425 0.6150 ;
        RECT 0.2850 0.1350 0.3450 0.1950 ;
        LAYER M1 ;
        RECT 1.2525 0.4500 1.2825 0.5700 ;
        RECT 1.1775 0.2550 1.2525 0.7650 ;
        RECT 1.0200 0.2550 1.1775 0.3300 ;
        RECT 1.0500 0.6900 1.1775 0.7650 ;
        RECT 0.9750 0.4050 1.1025 0.6150 ;
        RECT 0.9750 0.6900 1.0500 0.9000 ;
        RECT 0.9450 0.1500 1.0200 0.3300 ;
        RECT 0.9375 0.4050 0.9750 0.5400 ;
        RECT 0.6750 0.8250 0.9750 0.9000 ;
        RECT 0.6825 0.1500 0.9450 0.2550 ;
        RECT 0.7800 0.6375 0.9000 0.7500 ;
        RECT 0.7875 0.3600 0.8625 0.5625 ;
        RECT 0.6600 0.4875 0.7875 0.5625 ;
        RECT 0.6150 0.6750 0.7800 0.7500 ;
        RECT 0.6075 0.3300 0.6825 0.4125 ;
        RECT 0.5925 0.4875 0.6600 0.6000 ;
        RECT 0.5475 0.6750 0.6150 0.7650 ;
        RECT 0.5175 0.1500 0.6075 0.4125 ;
        RECT 0.4725 0.5250 0.5925 0.6000 ;
        RECT 0.1575 0.6900 0.5475 0.7650 ;
        RECT 0.4875 0.1500 0.5175 0.2250 ;
        RECT 0.2925 0.5250 0.4725 0.6150 ;
        RECT 0.3375 0.2850 0.4425 0.4050 ;
        RECT 0.1650 0.3300 0.3375 0.4050 ;
        RECT 0.1875 0.4800 0.2925 0.6150 ;
        RECT 0.1125 0.1500 0.1650 0.4050 ;
        RECT 0.1125 0.6900 0.1575 0.9000 ;
        RECT 0.0375 0.1500 0.1125 0.9000 ;
    END
END CKMUX2_1000


MACRO CKMUX2_1010
    CLASS CORE ;
    FOREIGN CKMUX2_1010 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.4700 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 1.3575 0.2025 1.4325 0.8325 ;
        RECT 1.3275 0.2025 1.3575 0.3825 ;
        RECT 1.3275 0.6675 1.3575 0.8325 ;
        END
    END Z
    PIN S
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.5025 0.5625 0.8625 0.6375 ;
        RECT 0.3975 0.4875 0.5025 0.6375 ;
        VIA 0.4500 0.5625 VIA12_square ;
        END
    END S
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.6525 0.4125 1.1175 0.4875 ;
        VIA 1.0200 0.4500 VIA12_square ;
        END
    END I1
    PIN I0
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.4275 0.2625 0.8925 0.3375 ;
        VIA 0.5625 0.3000 VIA12_square ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.2150 -0.0750 1.4700 0.0750 ;
        RECT 1.0950 -0.0750 1.2150 0.1800 ;
        RECT 0.3750 -0.0750 1.0950 0.0750 ;
        RECT 0.2550 -0.0750 0.3750 0.1800 ;
        RECT 0.0000 -0.0750 0.2550 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.2300 0.9750 1.4700 1.1250 ;
        RECT 1.1250 0.8400 1.2300 1.1250 ;
        RECT 0.3750 0.9750 1.1250 1.1250 ;
        RECT 0.2550 0.8625 0.3750 1.1250 ;
        RECT 0.0000 0.9750 0.2550 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.3350 0.2775 1.3950 0.3375 ;
        RECT 1.3350 0.7200 1.3950 0.7800 ;
        RECT 1.2225 0.4800 1.2825 0.5400 ;
        RECT 1.1250 0.1200 1.1850 0.1800 ;
        RECT 1.1250 0.8700 1.1850 0.9300 ;
        RECT 1.0200 0.4875 1.0800 0.5475 ;
        RECT 0.8100 0.6375 0.8700 0.6975 ;
        RECT 0.8025 0.3900 0.8625 0.4500 ;
        RECT 0.7050 0.1725 0.7650 0.2325 ;
        RECT 0.7050 0.8325 0.7650 0.8925 ;
        RECT 0.5925 0.3450 0.6525 0.4050 ;
        RECT 0.3825 0.3150 0.4425 0.3750 ;
        RECT 0.2850 0.8700 0.3450 0.9300 ;
        RECT 0.1875 0.5250 0.2475 0.5850 ;
        RECT 0.0750 0.1575 0.1350 0.2175 ;
        RECT 0.0750 0.7950 0.1350 0.8550 ;
        RECT 0.3825 0.5550 0.4425 0.6150 ;
        RECT 0.2850 0.1200 0.3450 0.1800 ;
        LAYER M1 ;
        RECT 1.2525 0.4500 1.2825 0.5700 ;
        RECT 1.1775 0.2550 1.2525 0.7650 ;
        RECT 1.0200 0.2550 1.1775 0.3300 ;
        RECT 1.0500 0.6900 1.1775 0.7650 ;
        RECT 0.9750 0.4050 1.1025 0.6150 ;
        RECT 0.9750 0.6900 1.0500 0.9000 ;
        RECT 0.9450 0.1500 1.0200 0.3300 ;
        RECT 0.9375 0.4050 0.9750 0.5400 ;
        RECT 0.6750 0.8250 0.9750 0.9000 ;
        RECT 0.6825 0.1500 0.9450 0.2550 ;
        RECT 0.7800 0.6375 0.9000 0.7500 ;
        RECT 0.7875 0.3600 0.8625 0.5625 ;
        RECT 0.6975 0.4875 0.7875 0.5625 ;
        RECT 0.6150 0.6750 0.7800 0.7500 ;
        RECT 0.6300 0.4875 0.6975 0.6000 ;
        RECT 0.6075 0.3300 0.6825 0.4125 ;
        RECT 0.4725 0.5250 0.6300 0.6000 ;
        RECT 0.5475 0.6750 0.6150 0.7650 ;
        RECT 0.5175 0.1500 0.6075 0.4125 ;
        RECT 0.1650 0.6900 0.5475 0.7650 ;
        RECT 0.4875 0.1500 0.5175 0.2250 ;
        RECT 0.2925 0.5250 0.4725 0.6150 ;
        RECT 0.3375 0.2850 0.4425 0.4050 ;
        RECT 0.1650 0.3300 0.3375 0.4050 ;
        RECT 0.1875 0.4800 0.2925 0.6150 ;
        RECT 0.1125 0.1500 0.1650 0.4050 ;
        RECT 0.1125 0.6900 0.1650 0.8625 ;
        RECT 0.0375 0.1500 0.1125 0.8625 ;
    END
END CKMUX2_1010


MACRO CKND2_0001
    CLASS CORE ;
    FOREIGN CKND2_0001 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.4700 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 0.5625 0.7125 1.0275 0.7875 ;
        RECT 0.4875 0.1575 0.5625 0.7875 ;
        RECT 0.3675 0.1575 0.4875 0.2325 ;
        VIA 0.5250 0.7050 VIA12_square ;
        VIA 0.4500 0.1950 VIA12_square ;
        END
    END ZN
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.3275 0.3675 1.4025 0.6825 ;
        RECT 0.7875 0.4875 1.3275 0.5925 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1500 0.4875 0.6825 0.5925 ;
        RECT 0.1425 0.3675 0.1500 0.5925 ;
        RECT 0.0675 0.3675 0.1425 0.6825 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.4025 -0.0750 1.4700 0.0750 ;
        RECT 1.3275 -0.0750 1.4025 0.2625 ;
        RECT 0.9975 -0.0750 1.3275 0.0750 ;
        RECT 0.8925 -0.0750 0.9975 0.2400 ;
        RECT 0.0000 -0.0750 0.8925 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.4025 0.9750 1.4700 1.1250 ;
        RECT 1.3275 0.7875 1.4025 1.1250 ;
        RECT 1.0050 0.9750 1.3275 1.1250 ;
        RECT 0.8850 0.8475 1.0050 1.1250 ;
        RECT 0.5850 0.9750 0.8850 1.1250 ;
        RECT 0.4650 0.8475 0.5850 1.1250 ;
        RECT 0.1425 0.9750 0.4650 1.1250 ;
        RECT 0.0675 0.7875 0.1425 1.1250 ;
        RECT 0.0000 0.9750 0.0675 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.3350 0.1725 1.3950 0.2325 ;
        RECT 1.3350 0.8175 1.3950 0.8775 ;
        RECT 1.2300 0.5100 1.2900 0.5700 ;
        RECT 1.1250 0.3300 1.1850 0.3900 ;
        RECT 1.1250 0.7725 1.1850 0.8325 ;
        RECT 1.0200 0.5100 1.0800 0.5700 ;
        RECT 0.9150 0.1575 0.9750 0.2175 ;
        RECT 0.9150 0.8550 0.9750 0.9150 ;
        RECT 0.8100 0.5100 0.8700 0.5700 ;
        RECT 0.7050 0.3300 0.7650 0.3900 ;
        RECT 0.7050 0.7725 0.7650 0.8325 ;
        RECT 0.6000 0.5100 0.6600 0.5700 ;
        RECT 0.4950 0.1650 0.5550 0.2250 ;
        RECT 0.4950 0.8550 0.5550 0.9150 ;
        RECT 0.3900 0.5100 0.4500 0.5700 ;
        RECT 0.2850 0.3300 0.3450 0.3900 ;
        RECT 0.2850 0.7725 0.3450 0.8325 ;
        RECT 0.1800 0.5100 0.2400 0.5700 ;
        RECT 0.0750 0.1800 0.1350 0.2400 ;
        RECT 0.0750 0.8175 0.1350 0.8775 ;
        LAYER M1 ;
        RECT 0.2550 0.3225 1.2150 0.3975 ;
        RECT 1.1025 0.6675 1.2075 0.8550 ;
        RECT 0.7875 0.6675 1.1025 0.7425 ;
        RECT 0.6825 0.6675 0.7875 0.8550 ;
        RECT 0.3675 0.6675 0.6825 0.7425 ;
        RECT 0.1575 0.1575 0.6075 0.2325 ;
        RECT 0.2625 0.6675 0.3675 0.8550 ;
        RECT 0.0525 0.1575 0.1575 0.2625 ;
    END
END CKND2_0001


MACRO CKND2_0011
    CLASS CORE ;
    FOREIGN CKND2_0011 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.0500 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.6975 0.6750 0.7725 0.8700 ;
        RECT 0.3675 0.6750 0.6975 0.7500 ;
        RECT 0.1125 0.3300 0.3750 0.4050 ;
        RECT 0.2625 0.6750 0.3675 0.8700 ;
        RECT 0.1125 0.6750 0.2625 0.7500 ;
        RECT 0.0375 0.3300 0.1125 0.7500 ;
        END
    END ZN
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.9075 0.4125 1.0125 0.6825 ;
        RECT 0.6000 0.4125 0.9075 0.5625 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.4950 0.2625 0.7575 0.3375 ;
        RECT 0.3900 0.2625 0.4950 0.6225 ;
        RECT 0.2925 0.2625 0.3900 0.3375 ;
        VIA 0.4425 0.5400 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.7950 -0.0750 1.0500 0.0750 ;
        RECT 0.6750 -0.0750 0.7950 0.1875 ;
        RECT 0.0000 -0.0750 0.6750 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.9825 0.9750 1.0500 1.1250 ;
        RECT 0.9075 0.8025 0.9825 1.1250 ;
        RECT 0.5850 0.9750 0.9075 1.1250 ;
        RECT 0.4650 0.8325 0.5850 1.1250 ;
        RECT 0.1650 0.9750 0.4650 1.1250 ;
        RECT 0.0450 0.8250 0.1650 1.1250 ;
        RECT 0.0000 0.9750 0.0450 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 0.9150 0.2100 0.9750 0.2700 ;
        RECT 0.9150 0.8325 0.9750 0.8925 ;
        RECT 0.8100 0.4650 0.8700 0.5250 ;
        RECT 0.7050 0.1200 0.7650 0.1800 ;
        RECT 0.7050 0.7800 0.7650 0.8400 ;
        RECT 0.6000 0.4650 0.6600 0.5250 ;
        RECT 0.4950 0.1575 0.5550 0.2175 ;
        RECT 0.4950 0.8400 0.5550 0.9000 ;
        RECT 0.3900 0.5100 0.4500 0.5700 ;
        RECT 0.2850 0.3300 0.3450 0.3900 ;
        RECT 0.2850 0.7800 0.3450 0.8400 ;
        RECT 0.1875 0.5100 0.2475 0.5700 ;
        RECT 0.0750 0.1725 0.1350 0.2325 ;
        RECT 0.0750 0.8325 0.1350 0.8925 ;
        LAYER M1 ;
        RECT 0.9075 0.1800 0.9825 0.3375 ;
        RECT 0.5850 0.2625 0.9075 0.3375 ;
        RECT 0.5100 0.1500 0.5850 0.3375 ;
        RECT 0.1875 0.4800 0.5250 0.6000 ;
        RECT 0.1650 0.1500 0.5100 0.2250 ;
        RECT 0.0450 0.1500 0.1650 0.2550 ;
    END
END CKND2_0011


MACRO CKND2_0100
    CLASS CORE ;
    FOREIGN CKND2_0100 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.5700 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 1.1025 0.3000 1.2600 0.4200 ;
        RECT 1.1025 0.6525 1.2600 0.7725 ;
        RECT 0.7875 0.3000 1.1025 0.7725 ;
        RECT 0.6300 0.3000 0.7875 0.4200 ;
        RECT 0.6300 0.6525 0.7875 0.7725 ;
        VIA 1.1025 0.3600 VIA12_slot ;
        VIA 1.1025 0.7125 VIA12_slot ;
        VIA 0.7875 0.3600 VIA12_slot ;
        VIA 0.7875 0.7125 VIA12_slot ;
        END
    END ZN
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 2.2050 0.5625 2.6700 0.6375 ;
        RECT 2.1000 0.4125 2.2050 0.6375 ;
        VIA 2.1525 0.4950 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1425 0.4950 1.7400 0.5700 ;
        RECT 0.0675 0.3675 0.1425 0.6825 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 3.3150 -0.0750 3.5700 0.0750 ;
        RECT 3.1950 -0.0750 3.3150 0.2250 ;
        RECT 2.8950 -0.0750 3.1950 0.0750 ;
        RECT 2.7750 -0.0750 2.8950 0.2250 ;
        RECT 2.4750 -0.0750 2.7750 0.0750 ;
        RECT 2.3550 -0.0750 2.4750 0.2250 ;
        RECT 2.0550 -0.0750 2.3550 0.0750 ;
        RECT 1.9350 -0.0750 2.0550 0.2250 ;
        RECT 0.0000 -0.0750 1.9350 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 3.5025 0.9750 3.5700 1.1250 ;
        RECT 3.4275 0.7875 3.5025 1.1250 ;
        RECT 3.1050 0.9750 3.4275 1.1250 ;
        RECT 2.9850 0.8475 3.1050 1.1250 ;
        RECT 2.6850 0.9750 2.9850 1.1250 ;
        RECT 2.5650 0.8475 2.6850 1.1250 ;
        RECT 2.2650 0.9750 2.5650 1.1250 ;
        RECT 2.1450 0.8475 2.2650 1.1250 ;
        RECT 1.8450 0.9750 2.1450 1.1250 ;
        RECT 1.7250 0.8475 1.8450 1.1250 ;
        RECT 1.4250 0.9750 1.7250 1.1250 ;
        RECT 1.3050 0.8475 1.4250 1.1250 ;
        RECT 1.0050 0.9750 1.3050 1.1250 ;
        RECT 0.8850 0.8475 1.0050 1.1250 ;
        RECT 0.5850 0.9750 0.8850 1.1250 ;
        RECT 0.4650 0.8475 0.5850 1.1250 ;
        RECT 0.1425 0.9750 0.4650 1.1250 ;
        RECT 0.0675 0.7875 0.1425 1.1250 ;
        RECT 0.0000 0.9750 0.0675 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 3.4350 0.2925 3.4950 0.3525 ;
        RECT 3.4350 0.8175 3.4950 0.8775 ;
        RECT 3.3300 0.4875 3.3900 0.5475 ;
        RECT 3.2250 0.1575 3.2850 0.2175 ;
        RECT 3.2250 0.7800 3.2850 0.8400 ;
        RECT 3.1200 0.4875 3.1800 0.5475 ;
        RECT 3.0150 0.3075 3.0750 0.3675 ;
        RECT 3.0150 0.8550 3.0750 0.9150 ;
        RECT 2.9100 0.4875 2.9700 0.5475 ;
        RECT 2.8050 0.1575 2.8650 0.2175 ;
        RECT 2.8050 0.7800 2.8650 0.8400 ;
        RECT 2.7000 0.4875 2.7600 0.5475 ;
        RECT 2.5950 0.3075 2.6550 0.3675 ;
        RECT 2.5950 0.8550 2.6550 0.9150 ;
        RECT 2.4900 0.4875 2.5500 0.5475 ;
        RECT 2.3850 0.1575 2.4450 0.2175 ;
        RECT 2.3850 0.7800 2.4450 0.8400 ;
        RECT 2.2800 0.4875 2.3400 0.5475 ;
        RECT 2.1750 0.3075 2.2350 0.3675 ;
        RECT 2.1750 0.8550 2.2350 0.9150 ;
        RECT 2.0700 0.4875 2.1300 0.5475 ;
        RECT 1.9650 0.1575 2.0250 0.2175 ;
        RECT 1.9650 0.7800 2.0250 0.8400 ;
        RECT 1.8600 0.4875 1.9200 0.5475 ;
        RECT 1.7550 0.2325 1.8150 0.2925 ;
        RECT 1.7550 0.8550 1.8150 0.9150 ;
        RECT 1.6500 0.5025 1.7100 0.5625 ;
        RECT 1.5450 0.3300 1.6050 0.3900 ;
        RECT 1.5450 0.7950 1.6050 0.8550 ;
        RECT 1.4400 0.5025 1.5000 0.5625 ;
        RECT 1.3350 0.1575 1.3950 0.2175 ;
        RECT 1.3350 0.8550 1.3950 0.9150 ;
        RECT 1.2300 0.5025 1.2900 0.5625 ;
        RECT 1.1250 0.3300 1.1850 0.3900 ;
        RECT 1.1250 0.7950 1.1850 0.8550 ;
        RECT 1.0200 0.5025 1.0800 0.5625 ;
        RECT 0.9150 0.1575 0.9750 0.2175 ;
        RECT 0.9150 0.8550 0.9750 0.9150 ;
        RECT 0.8100 0.5025 0.8700 0.5625 ;
        RECT 0.7050 0.3300 0.7650 0.3900 ;
        RECT 0.7050 0.7950 0.7650 0.8550 ;
        RECT 0.0750 0.1725 0.1350 0.2325 ;
        RECT 0.0750 0.8250 0.1350 0.8850 ;
        RECT 0.6000 0.5025 0.6600 0.5625 ;
        RECT 0.4950 0.1575 0.5550 0.2175 ;
        RECT 0.4950 0.8550 0.5550 0.9150 ;
        RECT 0.3900 0.5025 0.4500 0.5625 ;
        RECT 0.2850 0.3300 0.3450 0.3900 ;
        RECT 0.2850 0.7950 0.3450 0.8550 ;
        RECT 0.1800 0.5025 0.2400 0.5625 ;
        LAYER M1 ;
        RECT 3.4125 0.2700 3.5175 0.3750 ;
        RECT 1.8225 0.3000 3.4125 0.3750 ;
        RECT 1.8525 0.4575 3.4050 0.5775 ;
        RECT 3.2025 0.6525 3.3075 0.8625 ;
        RECT 2.8875 0.6525 3.2025 0.7725 ;
        RECT 2.7825 0.6525 2.8875 0.8625 ;
        RECT 2.4675 0.6525 2.7825 0.7725 ;
        RECT 2.3625 0.6525 2.4675 0.8625 ;
        RECT 2.0475 0.6525 2.3625 0.7725 ;
        RECT 1.9425 0.6525 2.0475 0.8625 ;
        RECT 1.6275 0.6525 1.9425 0.7725 ;
        RECT 1.7475 0.1500 1.8225 0.3750 ;
        RECT 0.1575 0.1500 1.7475 0.2250 ;
        RECT 0.2550 0.3000 1.6350 0.4200 ;
        RECT 1.5225 0.6525 1.6275 0.8775 ;
        RECT 1.2075 0.6525 1.5225 0.7725 ;
        RECT 1.1025 0.6525 1.2075 0.8775 ;
        RECT 0.7875 0.6525 1.1025 0.7725 ;
        RECT 0.6825 0.6525 0.7875 0.8775 ;
        RECT 0.3675 0.6525 0.6825 0.7725 ;
        RECT 0.2625 0.6525 0.3675 0.8775 ;
        RECT 0.0525 0.1500 0.1575 0.2550 ;
        LAYER M2 ;
        RECT 1.1325 0.3000 1.2600 0.4200 ;
        RECT 1.1325 0.6525 1.2600 0.7725 ;
        RECT 0.6300 0.3000 0.7575 0.4200 ;
        RECT 0.6300 0.6525 0.7575 0.7725 ;
    END
END CKND2_0100


MACRO CKND2_0111
    CLASS CORE ;
    FOREIGN CKND2_0111 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.8900 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 1.2075 0.2700 1.5225 0.7950 ;
        VIA 1.3650 0.3525 VIA12_slot ;
        VIA 1.3650 0.7125 VIA12_slot ;
        END
    END ZN
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.4725 0.4125 0.9225 0.4875 ;
        RECT 0.3675 0.4125 0.4725 0.6225 ;
        VIA 0.4200 0.5400 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.7475 0.3675 1.8225 0.6825 ;
        RECT 0.9975 0.4800 1.7475 0.5850 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.7950 -0.0750 1.8900 0.0750 ;
        RECT 0.6750 -0.0750 0.7950 0.2250 ;
        RECT 0.3750 -0.0750 0.6750 0.0750 ;
        RECT 0.2550 -0.0750 0.3750 0.2250 ;
        RECT 0.0000 -0.0750 0.2550 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.8225 0.9750 1.8900 1.1250 ;
        RECT 1.7475 0.8025 1.8225 1.1250 ;
        RECT 1.4250 0.9750 1.7475 1.1250 ;
        RECT 1.3050 0.8475 1.4250 1.1250 ;
        RECT 1.0050 0.9750 1.3050 1.1250 ;
        RECT 0.8850 0.8400 1.0050 1.1250 ;
        RECT 0.5850 0.9750 0.8850 1.1250 ;
        RECT 0.4650 0.8400 0.5850 1.1250 ;
        RECT 0.1425 0.9750 0.4650 1.1250 ;
        RECT 0.0675 0.8025 0.1425 1.1250 ;
        RECT 0.0000 0.9750 0.0675 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.7550 0.1725 1.8150 0.2325 ;
        RECT 1.7550 0.8325 1.8150 0.8925 ;
        RECT 1.6500 0.5025 1.7100 0.5625 ;
        RECT 1.5450 0.3225 1.6050 0.3825 ;
        RECT 1.5450 0.7800 1.6050 0.8400 ;
        RECT 1.4400 0.5025 1.5000 0.5625 ;
        RECT 1.3350 0.1575 1.3950 0.2175 ;
        RECT 1.3350 0.8550 1.3950 0.9150 ;
        RECT 1.2300 0.5025 1.2900 0.5625 ;
        RECT 1.1250 0.3225 1.1850 0.3825 ;
        RECT 1.1250 0.7800 1.1850 0.8400 ;
        RECT 1.0200 0.5025 1.0800 0.5625 ;
        RECT 0.9150 0.2325 0.9750 0.2925 ;
        RECT 0.9150 0.8475 0.9750 0.9075 ;
        RECT 0.8100 0.5025 0.8700 0.5625 ;
        RECT 0.7050 0.1575 0.7650 0.2175 ;
        RECT 0.7050 0.7800 0.7650 0.8400 ;
        RECT 0.6000 0.5025 0.6600 0.5625 ;
        RECT 0.4950 0.3075 0.5550 0.3675 ;
        RECT 0.4950 0.8475 0.5550 0.9075 ;
        RECT 0.3900 0.5025 0.4500 0.5625 ;
        RECT 0.2850 0.1575 0.3450 0.2175 ;
        RECT 0.2850 0.7800 0.3450 0.8400 ;
        RECT 0.1800 0.5025 0.2400 0.5625 ;
        RECT 0.0750 0.2925 0.1350 0.3525 ;
        RECT 0.0750 0.8325 0.1350 0.8925 ;
        LAYER M1 ;
        RECT 1.7325 0.1500 1.8375 0.2550 ;
        RECT 0.9825 0.1500 1.7325 0.2250 ;
        RECT 1.1025 0.3000 1.6275 0.4050 ;
        RECT 1.5225 0.6600 1.6275 0.8625 ;
        RECT 1.2075 0.6600 1.5225 0.7650 ;
        RECT 1.1025 0.6600 1.2075 0.8625 ;
        RECT 0.7875 0.6600 1.1025 0.7650 ;
        RECT 0.9075 0.1500 0.9825 0.3750 ;
        RECT 0.1575 0.3000 0.9075 0.3750 ;
        RECT 0.1500 0.4800 0.8925 0.5850 ;
        RECT 0.6825 0.6600 0.7875 0.8625 ;
        RECT 0.3675 0.6600 0.6825 0.7650 ;
        RECT 0.2625 0.6600 0.3675 0.8625 ;
        RECT 0.0525 0.2700 0.1575 0.3750 ;
    END
END CKND2_0111


MACRO CKND2_1000
    CLASS CORE ;
    FOREIGN CKND2_1000 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.6300 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.5175 0.1725 0.5925 0.7425 ;
        RECT 0.4875 0.1725 0.5175 0.3825 ;
        RECT 0.3675 0.6675 0.5175 0.7425 ;
        RECT 0.2625 0.6675 0.3675 0.8925 ;
        END
    END ZN
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1425 0.4575 0.2325 0.5925 ;
        RECT 0.0675 0.3675 0.1425 0.6825 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.3825 0.4425 0.4425 0.5925 ;
        RECT 0.3075 0.2175 0.3825 0.5925 ;
        RECT 0.2775 0.2175 0.3075 0.3825 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.1425 -0.0750 0.6300 0.0750 ;
        RECT 0.0675 -0.0750 0.1425 0.2475 ;
        RECT 0.0000 -0.0750 0.0675 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.5925 0.9750 0.6300 1.1250 ;
        RECT 0.4575 0.8175 0.5925 1.1250 ;
        RECT 0.1425 0.9750 0.4575 1.1250 ;
        RECT 0.0675 0.8025 0.1425 1.1250 ;
        RECT 0.0000 0.9750 0.0675 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 0.4950 0.2025 0.5550 0.2625 ;
        RECT 0.4950 0.8325 0.5550 0.8925 ;
        RECT 0.3825 0.4875 0.4425 0.5475 ;
        RECT 0.2850 0.8025 0.3450 0.8625 ;
        RECT 0.1725 0.4875 0.2325 0.5475 ;
        RECT 0.0750 0.1575 0.1350 0.2175 ;
        RECT 0.0750 0.8325 0.1350 0.8925 ;
    END
END CKND2_1000


MACRO CKND2_1010
    CLASS CORE ;
    FOREIGN CKND2_1010 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.6300 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.5175 0.1800 0.5925 0.7425 ;
        RECT 0.4875 0.1800 0.5175 0.3825 ;
        RECT 0.3525 0.6675 0.5175 0.7425 ;
        RECT 0.2775 0.6675 0.3525 0.8700 ;
        END
    END ZN
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1425 0.4575 0.2325 0.5925 ;
        RECT 0.0675 0.3675 0.1425 0.6825 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.3825 0.4425 0.4425 0.5925 ;
        RECT 0.3075 0.2175 0.3825 0.5925 ;
        RECT 0.2775 0.2175 0.3075 0.3825 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.1425 -0.0750 0.6300 0.0750 ;
        RECT 0.0675 -0.0750 0.1425 0.2475 ;
        RECT 0.0000 -0.0750 0.0675 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.5925 0.9750 0.6300 1.1250 ;
        RECT 0.4575 0.8175 0.5925 1.1250 ;
        RECT 0.1425 0.9750 0.4575 1.1250 ;
        RECT 0.0675 0.8025 0.1425 1.1250 ;
        RECT 0.0000 0.9750 0.0675 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 0.4950 0.2100 0.5550 0.2700 ;
        RECT 0.4950 0.8325 0.5550 0.8925 ;
        RECT 0.3825 0.4875 0.4425 0.5475 ;
        RECT 0.2850 0.7650 0.3450 0.8250 ;
        RECT 0.1725 0.4875 0.2325 0.5475 ;
        RECT 0.0750 0.1575 0.1350 0.2175 ;
        RECT 0.0750 0.8325 0.1350 0.8925 ;
    END
END CKND2_1010


MACRO CKN_0000
    CLASS CORE ;
    FOREIGN CKN_0000 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.4100 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 2.3625 0.2775 2.5200 0.3975 ;
        RECT 2.3625 0.6525 2.5200 0.7725 ;
        RECT 2.0475 0.2775 2.3625 0.7725 ;
        RECT 1.8900 0.2775 2.0475 0.3975 ;
        RECT 1.8900 0.6525 2.0475 0.7725 ;
        VIA 2.3625 0.3375 VIA12_slot ;
        VIA 2.3625 0.7125 VIA12_slot ;
        VIA 2.0475 0.3375 VIA12_slot ;
        VIA 2.0475 0.7125 VIA12_slot ;
        END
    END ZN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1425 0.4725 4.3050 0.5475 ;
        RECT 0.0675 0.3675 0.1425 0.6825 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 4.3650 -0.0750 4.4100 0.0750 ;
        RECT 4.2450 -0.0750 4.3650 0.2925 ;
        RECT 3.9450 -0.0750 4.2450 0.0750 ;
        RECT 3.8250 -0.0750 3.9450 0.2025 ;
        RECT 3.5250 -0.0750 3.8250 0.0750 ;
        RECT 3.4050 -0.0750 3.5250 0.2025 ;
        RECT 3.1050 -0.0750 3.4050 0.0750 ;
        RECT 2.9850 -0.0750 3.1050 0.2025 ;
        RECT 2.6850 -0.0750 2.9850 0.0750 ;
        RECT 2.5650 -0.0750 2.6850 0.2025 ;
        RECT 2.2650 -0.0750 2.5650 0.0750 ;
        RECT 2.1450 -0.0750 2.2650 0.2025 ;
        RECT 1.8450 -0.0750 2.1450 0.0750 ;
        RECT 1.7250 -0.0750 1.8450 0.2025 ;
        RECT 1.4250 -0.0750 1.7250 0.0750 ;
        RECT 1.3050 -0.0750 1.4250 0.2025 ;
        RECT 1.0050 -0.0750 1.3050 0.0750 ;
        RECT 0.8850 -0.0750 1.0050 0.2025 ;
        RECT 0.5850 -0.0750 0.8850 0.0750 ;
        RECT 0.4650 -0.0750 0.5850 0.2025 ;
        RECT 0.1425 -0.0750 0.4650 0.0750 ;
        RECT 0.0675 -0.0750 0.1425 0.2475 ;
        RECT 0.0000 -0.0750 0.0675 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 4.3650 0.9750 4.4100 1.1250 ;
        RECT 4.2450 0.6600 4.3650 1.1250 ;
        RECT 3.9450 0.9750 4.2450 1.1250 ;
        RECT 3.8250 0.8475 3.9450 1.1250 ;
        RECT 3.5250 0.9750 3.8250 1.1250 ;
        RECT 3.4050 0.8475 3.5250 1.1250 ;
        RECT 3.1050 0.9750 3.4050 1.1250 ;
        RECT 2.9850 0.8475 3.1050 1.1250 ;
        RECT 2.6850 0.9750 2.9850 1.1250 ;
        RECT 2.5650 0.8475 2.6850 1.1250 ;
        RECT 2.2650 0.9750 2.5650 1.1250 ;
        RECT 2.1450 0.8475 2.2650 1.1250 ;
        RECT 1.8450 0.9750 2.1450 1.1250 ;
        RECT 1.7250 0.8475 1.8450 1.1250 ;
        RECT 1.4250 0.9750 1.7250 1.1250 ;
        RECT 1.3050 0.8475 1.4250 1.1250 ;
        RECT 1.0050 0.9750 1.3050 1.1250 ;
        RECT 0.8850 0.8475 1.0050 1.1250 ;
        RECT 0.5850 0.9750 0.8850 1.1250 ;
        RECT 0.4650 0.8475 0.5850 1.1250 ;
        RECT 0.1425 0.9750 0.4650 1.1250 ;
        RECT 0.0675 0.8025 0.1425 1.1250 ;
        RECT 0.0000 0.9750 0.0675 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 4.2750 0.2250 4.3350 0.2850 ;
        RECT 4.2750 0.6675 4.3350 0.7275 ;
        RECT 4.2750 0.8325 4.3350 0.8925 ;
        RECT 4.1700 0.4800 4.2300 0.5400 ;
        RECT 4.0650 0.3075 4.1250 0.3675 ;
        RECT 4.0650 0.6825 4.1250 0.7425 ;
        RECT 3.9600 0.4800 4.0200 0.5400 ;
        RECT 3.8550 0.1350 3.9150 0.1950 ;
        RECT 3.8550 0.8550 3.9150 0.9150 ;
        RECT 3.7500 0.4800 3.8100 0.5400 ;
        RECT 3.6450 0.3075 3.7050 0.3675 ;
        RECT 3.6450 0.6825 3.7050 0.7425 ;
        RECT 3.5400 0.4800 3.6000 0.5400 ;
        RECT 3.4350 0.1350 3.4950 0.1950 ;
        RECT 3.4350 0.8550 3.4950 0.9150 ;
        RECT 3.3300 0.4800 3.3900 0.5400 ;
        RECT 3.2250 0.3075 3.2850 0.3675 ;
        RECT 3.2250 0.6825 3.2850 0.7425 ;
        RECT 3.1200 0.4800 3.1800 0.5400 ;
        RECT 3.0150 0.1350 3.0750 0.1950 ;
        RECT 3.0150 0.8550 3.0750 0.9150 ;
        RECT 2.9100 0.4800 2.9700 0.5400 ;
        RECT 2.8050 0.3075 2.8650 0.3675 ;
        RECT 2.8050 0.6825 2.8650 0.7425 ;
        RECT 2.7000 0.4800 2.7600 0.5400 ;
        RECT 2.5950 0.1350 2.6550 0.1950 ;
        RECT 2.5950 0.8550 2.6550 0.9150 ;
        RECT 2.4900 0.4800 2.5500 0.5400 ;
        RECT 2.3850 0.3075 2.4450 0.3675 ;
        RECT 2.3850 0.6825 2.4450 0.7425 ;
        RECT 2.2800 0.4800 2.3400 0.5400 ;
        RECT 2.1750 0.1350 2.2350 0.1950 ;
        RECT 2.1750 0.8550 2.2350 0.9150 ;
        RECT 2.0700 0.4800 2.1300 0.5400 ;
        RECT 1.9650 0.3075 2.0250 0.3675 ;
        RECT 1.9650 0.6825 2.0250 0.7425 ;
        RECT 1.8600 0.4800 1.9200 0.5400 ;
        RECT 1.7550 0.1350 1.8150 0.1950 ;
        RECT 1.7550 0.8550 1.8150 0.9150 ;
        RECT 1.6500 0.4800 1.7100 0.5400 ;
        RECT 1.5450 0.3075 1.6050 0.3675 ;
        RECT 1.5450 0.6825 1.6050 0.7425 ;
        RECT 1.4400 0.4800 1.5000 0.5400 ;
        RECT 1.3350 0.1350 1.3950 0.1950 ;
        RECT 1.3350 0.8550 1.3950 0.9150 ;
        RECT 1.2300 0.4800 1.2900 0.5400 ;
        RECT 1.1250 0.3075 1.1850 0.3675 ;
        RECT 1.1250 0.6825 1.1850 0.7425 ;
        RECT 1.0200 0.4800 1.0800 0.5400 ;
        RECT 0.9150 0.1350 0.9750 0.1950 ;
        RECT 0.9150 0.8550 0.9750 0.9150 ;
        RECT 0.8100 0.4800 0.8700 0.5400 ;
        RECT 0.7050 0.3075 0.7650 0.3675 ;
        RECT 0.7050 0.6825 0.7650 0.7425 ;
        RECT 0.6000 0.4800 0.6600 0.5400 ;
        RECT 0.4950 0.1350 0.5550 0.1950 ;
        RECT 0.4950 0.8550 0.5550 0.9150 ;
        RECT 0.3900 0.4800 0.4500 0.5400 ;
        RECT 0.2850 0.3075 0.3450 0.3675 ;
        RECT 0.2850 0.6825 0.3450 0.7425 ;
        RECT 0.1800 0.4800 0.2400 0.5400 ;
        RECT 0.0750 0.1575 0.1350 0.2175 ;
        RECT 0.0750 0.8325 0.1350 0.8925 ;
        LAYER M1 ;
        RECT 0.2775 0.2775 4.1400 0.3975 ;
        RECT 0.2775 0.6525 4.1400 0.7725 ;
        LAYER M2 ;
        RECT 2.3925 0.2775 2.5200 0.3975 ;
        RECT 2.3925 0.6525 2.5200 0.7725 ;
        RECT 1.8900 0.2775 2.0175 0.3975 ;
        RECT 1.8900 0.6525 2.0175 0.7725 ;
    END
END CKN_0000


MACRO CKN_0001
    CLASS CORE ;
    FOREIGN CKN_0001 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.8400 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.7725 0.2100 0.8025 0.7275 ;
        RECT 0.7275 0.2100 0.7725 0.8325 ;
        RECT 0.6750 0.2100 0.7275 0.3750 ;
        RECT 0.6975 0.6525 0.7275 0.8325 ;
        RECT 0.3525 0.6525 0.6975 0.7275 ;
        RECT 0.3525 0.3000 0.6750 0.3750 ;
        RECT 0.2775 0.1875 0.3525 0.3750 ;
        RECT 0.2775 0.6525 0.3525 0.8325 ;
        END
    END ZN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1425 0.4575 0.6525 0.5775 ;
        RECT 0.0675 0.3675 0.1425 0.6825 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.5850 -0.0750 0.8400 0.0750 ;
        RECT 0.4650 -0.0750 0.5850 0.2250 ;
        RECT 0.1425 -0.0750 0.4650 0.0750 ;
        RECT 0.0675 -0.0750 0.1425 0.2475 ;
        RECT 0.0000 -0.0750 0.0675 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.5775 0.9750 0.8400 1.1250 ;
        RECT 0.4725 0.8025 0.5775 1.1250 ;
        RECT 0.1425 0.9750 0.4725 1.1250 ;
        RECT 0.0675 0.8025 0.1425 1.1250 ;
        RECT 0.0000 0.9750 0.0675 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 0.7050 0.2175 0.7650 0.2775 ;
        RECT 0.7050 0.7425 0.7650 0.8025 ;
        RECT 0.5925 0.4875 0.6525 0.5475 ;
        RECT 0.4950 0.1575 0.5550 0.2175 ;
        RECT 0.4950 0.8250 0.5550 0.8850 ;
        RECT 0.3900 0.4875 0.4500 0.5475 ;
        RECT 0.2850 0.2250 0.3450 0.2850 ;
        RECT 0.2850 0.7425 0.3450 0.8025 ;
        RECT 0.1800 0.4875 0.2400 0.5475 ;
        RECT 0.0750 0.1575 0.1350 0.2175 ;
        RECT 0.0750 0.8325 0.1350 0.8925 ;
    END
END CKN_0001


MACRO CKN_0011
    CLASS CORE ;
    FOREIGN CKN_0011 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.6300 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.5175 0.3075 0.5925 0.7275 ;
        RECT 0.3525 0.3075 0.5175 0.3825 ;
        RECT 0.3525 0.6525 0.5175 0.7275 ;
        RECT 0.2775 0.1875 0.3525 0.3825 ;
        RECT 0.2775 0.6525 0.3525 0.8325 ;
        END
    END ZN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1425 0.4575 0.4425 0.5775 ;
        RECT 0.0675 0.3675 0.1425 0.6825 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.5850 -0.0750 0.6300 0.0750 ;
        RECT 0.4650 -0.0750 0.5850 0.2325 ;
        RECT 0.1425 -0.0750 0.4650 0.0750 ;
        RECT 0.0675 -0.0750 0.1425 0.2475 ;
        RECT 0.0000 -0.0750 0.0675 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.5775 0.9750 0.6300 1.1250 ;
        RECT 0.4725 0.8025 0.5775 1.1250 ;
        RECT 0.1425 0.9750 0.4725 1.1250 ;
        RECT 0.0675 0.8025 0.1425 1.1250 ;
        RECT 0.0000 0.9750 0.0675 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 0.4950 0.1575 0.5550 0.2175 ;
        RECT 0.4950 0.8250 0.5550 0.8850 ;
        RECT 0.3825 0.4875 0.4425 0.5475 ;
        RECT 0.2850 0.2250 0.3450 0.2850 ;
        RECT 0.2850 0.7425 0.3450 0.8025 ;
        RECT 0.1800 0.4875 0.2400 0.5475 ;
        RECT 0.0750 0.1575 0.1350 0.2175 ;
        RECT 0.0750 0.8325 0.1350 0.8925 ;
    END
END CKN_0011


MACRO CKN_0100
    CLASS CORE ;
    FOREIGN CKN_0100 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.8900 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 1.1025 0.2775 1.2600 0.3975 ;
        RECT 1.1025 0.6525 1.2600 0.7725 ;
        RECT 0.7875 0.2775 1.1025 0.7725 ;
        RECT 0.6300 0.2775 0.7875 0.3975 ;
        RECT 0.6300 0.6525 0.7875 0.7725 ;
        VIA 1.1025 0.3375 VIA12_slot ;
        VIA 1.1025 0.7125 VIA12_slot ;
        VIA 0.7875 0.3375 VIA12_slot ;
        VIA 0.7875 0.7125 VIA12_slot ;
        END
    END ZN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1425 0.4725 1.7850 0.5475 ;
        RECT 0.0675 0.3675 0.1425 0.6825 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.8450 -0.0750 1.8900 0.0750 ;
        RECT 1.7250 -0.0750 1.8450 0.2925 ;
        RECT 1.4250 -0.0750 1.7250 0.0750 ;
        RECT 1.3050 -0.0750 1.4250 0.2025 ;
        RECT 1.0050 -0.0750 1.3050 0.0750 ;
        RECT 0.8850 -0.0750 1.0050 0.2025 ;
        RECT 0.5850 -0.0750 0.8850 0.0750 ;
        RECT 0.4650 -0.0750 0.5850 0.2025 ;
        RECT 0.1425 -0.0750 0.4650 0.0750 ;
        RECT 0.0675 -0.0750 0.1425 0.2475 ;
        RECT 0.0000 -0.0750 0.0675 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.8450 0.9750 1.8900 1.1250 ;
        RECT 1.7250 0.6600 1.8450 1.1250 ;
        RECT 1.4250 0.9750 1.7250 1.1250 ;
        RECT 1.3050 0.8475 1.4250 1.1250 ;
        RECT 1.0050 0.9750 1.3050 1.1250 ;
        RECT 0.8850 0.8475 1.0050 1.1250 ;
        RECT 0.5850 0.9750 0.8850 1.1250 ;
        RECT 0.4650 0.8475 0.5850 1.1250 ;
        RECT 0.1425 0.9750 0.4650 1.1250 ;
        RECT 0.0675 0.8025 0.1425 1.1250 ;
        RECT 0.0000 0.9750 0.0675 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.7550 0.2250 1.8150 0.2850 ;
        RECT 1.7550 0.6675 1.8150 0.7275 ;
        RECT 1.7550 0.8325 1.8150 0.8925 ;
        RECT 1.6500 0.4800 1.7100 0.5400 ;
        RECT 1.5450 0.2625 1.6050 0.3225 ;
        RECT 1.5450 0.6825 1.6050 0.7425 ;
        RECT 1.4400 0.4800 1.5000 0.5400 ;
        RECT 1.3350 0.1350 1.3950 0.1950 ;
        RECT 1.3350 0.8550 1.3950 0.9150 ;
        RECT 1.2300 0.4800 1.2900 0.5400 ;
        RECT 1.1250 0.2625 1.1850 0.3225 ;
        RECT 1.1250 0.6825 1.1850 0.7425 ;
        RECT 1.0200 0.4800 1.0800 0.5400 ;
        RECT 0.9150 0.1350 0.9750 0.1950 ;
        RECT 0.9150 0.8550 0.9750 0.9150 ;
        RECT 0.8100 0.4800 0.8700 0.5400 ;
        RECT 0.7050 0.2625 0.7650 0.3225 ;
        RECT 0.7050 0.6825 0.7650 0.7425 ;
        RECT 0.6000 0.4800 0.6600 0.5400 ;
        RECT 0.4950 0.1350 0.5550 0.1950 ;
        RECT 0.4950 0.8550 0.5550 0.9150 ;
        RECT 0.3900 0.4800 0.4500 0.5400 ;
        RECT 0.2850 0.2625 0.3450 0.3225 ;
        RECT 0.2850 0.6825 0.3450 0.7425 ;
        RECT 0.1800 0.4800 0.2400 0.5400 ;
        RECT 0.0750 0.1575 0.1350 0.2175 ;
        RECT 0.0750 0.8325 0.1350 0.8925 ;
        LAYER M1 ;
        RECT 1.5150 0.2325 1.6350 0.3975 ;
        RECT 0.2775 0.6525 1.6200 0.7725 ;
        RECT 0.3750 0.2775 0.6750 0.3975 ;
        RECT 0.2550 0.2325 0.3750 0.3975 ;
        RECT 1.2150 0.2775 1.5150 0.3975 ;
        RECT 1.0950 0.2325 1.2150 0.3975 ;
        RECT 0.7950 0.2775 1.0950 0.3975 ;
        RECT 0.6750 0.2325 0.7950 0.3975 ;
        LAYER M2 ;
        RECT 1.1325 0.2775 1.2600 0.3975 ;
        RECT 1.1325 0.6525 1.2600 0.7725 ;
        RECT 0.6300 0.2775 0.7575 0.3975 ;
        RECT 0.6300 0.6525 0.7575 0.7725 ;
    END
END CKN_0100


MACRO CKN_0101
    CLASS CORE ;
    FOREIGN CKN_0101 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.7300 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 1.5225 0.2775 1.6800 0.3975 ;
        RECT 1.5225 0.6525 1.6800 0.7725 ;
        RECT 1.2075 0.2775 1.5225 0.7725 ;
        RECT 1.0500 0.2775 1.2075 0.3975 ;
        RECT 1.0500 0.6525 1.2075 0.7725 ;
        VIA 1.5225 0.3375 VIA12_slot ;
        VIA 1.5225 0.7125 VIA12_slot ;
        VIA 1.2075 0.3375 VIA12_slot ;
        VIA 1.2075 0.7125 VIA12_slot ;
        END
    END ZN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1425 0.4725 2.6250 0.5475 ;
        RECT 0.0675 0.3675 0.1425 0.6825 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 2.6850 -0.0750 2.7300 0.0750 ;
        RECT 2.5650 -0.0750 2.6850 0.2925 ;
        RECT 2.2650 -0.0750 2.5650 0.0750 ;
        RECT 2.1450 -0.0750 2.2650 0.2025 ;
        RECT 1.8450 -0.0750 2.1450 0.0750 ;
        RECT 1.7250 -0.0750 1.8450 0.2025 ;
        RECT 1.4250 -0.0750 1.7250 0.0750 ;
        RECT 1.3050 -0.0750 1.4250 0.2025 ;
        RECT 1.0050 -0.0750 1.3050 0.0750 ;
        RECT 0.8850 -0.0750 1.0050 0.2025 ;
        RECT 0.5850 -0.0750 0.8850 0.0750 ;
        RECT 0.4650 -0.0750 0.5850 0.2025 ;
        RECT 0.1425 -0.0750 0.4650 0.0750 ;
        RECT 0.0675 -0.0750 0.1425 0.2475 ;
        RECT 0.0000 -0.0750 0.0675 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 2.6850 0.9750 2.7300 1.1250 ;
        RECT 2.5650 0.6600 2.6850 1.1250 ;
        RECT 2.2650 0.9750 2.5650 1.1250 ;
        RECT 2.1450 0.8475 2.2650 1.1250 ;
        RECT 1.8450 0.9750 2.1450 1.1250 ;
        RECT 1.7250 0.8475 1.8450 1.1250 ;
        RECT 1.4250 0.9750 1.7250 1.1250 ;
        RECT 1.3050 0.8475 1.4250 1.1250 ;
        RECT 1.0050 0.9750 1.3050 1.1250 ;
        RECT 0.8850 0.8475 1.0050 1.1250 ;
        RECT 0.5850 0.9750 0.8850 1.1250 ;
        RECT 0.4650 0.8475 0.5850 1.1250 ;
        RECT 0.1425 0.9750 0.4650 1.1250 ;
        RECT 0.0675 0.8025 0.1425 1.1250 ;
        RECT 0.0000 0.9750 0.0675 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 2.5950 0.2175 2.6550 0.2775 ;
        RECT 2.5950 0.6675 2.6550 0.7275 ;
        RECT 2.5950 0.8325 2.6550 0.8925 ;
        RECT 2.3850 0.6825 2.4450 0.7425 ;
        RECT 2.2800 0.4800 2.3400 0.5400 ;
        RECT 2.1750 0.1350 2.2350 0.1950 ;
        RECT 2.1750 0.8550 2.2350 0.9150 ;
        RECT 2.0700 0.4800 2.1300 0.5400 ;
        RECT 1.9650 0.3075 2.0250 0.3675 ;
        RECT 1.9650 0.6825 2.0250 0.7425 ;
        RECT 1.8600 0.4800 1.9200 0.5400 ;
        RECT 1.7550 0.1350 1.8150 0.1950 ;
        RECT 1.7550 0.8550 1.8150 0.9150 ;
        RECT 1.6500 0.4800 1.7100 0.5400 ;
        RECT 1.5450 0.3075 1.6050 0.3675 ;
        RECT 1.5450 0.6825 1.6050 0.7425 ;
        RECT 1.4400 0.4800 1.5000 0.5400 ;
        RECT 1.3350 0.1350 1.3950 0.1950 ;
        RECT 1.3350 0.8550 1.3950 0.9150 ;
        RECT 1.2300 0.4800 1.2900 0.5400 ;
        RECT 1.1250 0.3075 1.1850 0.3675 ;
        RECT 1.1250 0.6825 1.1850 0.7425 ;
        RECT 1.0200 0.4800 1.0800 0.5400 ;
        RECT 0.9150 0.1350 0.9750 0.1950 ;
        RECT 0.9150 0.8550 0.9750 0.9150 ;
        RECT 0.8100 0.4800 0.8700 0.5400 ;
        RECT 0.7050 0.3075 0.7650 0.3675 ;
        RECT 0.7050 0.6825 0.7650 0.7425 ;
        RECT 0.6000 0.4800 0.6600 0.5400 ;
        RECT 0.4950 0.1350 0.5550 0.1950 ;
        RECT 0.4950 0.8550 0.5550 0.9150 ;
        RECT 0.3900 0.4800 0.4500 0.5400 ;
        RECT 0.2850 0.3075 0.3450 0.3675 ;
        RECT 0.2850 0.6825 0.3450 0.7425 ;
        RECT 0.1800 0.4800 0.2400 0.5400 ;
        RECT 0.0750 0.1575 0.1350 0.2175 ;
        RECT 0.0750 0.8325 0.1350 0.8925 ;
        RECT 2.4900 0.4800 2.5500 0.5400 ;
        RECT 2.3850 0.3075 2.4450 0.3675 ;
        LAYER M1 ;
        RECT 0.2775 0.2775 2.4600 0.3975 ;
        RECT 0.2775 0.6525 2.4600 0.7725 ;
        LAYER M2 ;
        RECT 1.5525 0.2775 1.6800 0.3975 ;
        RECT 1.5525 0.6525 1.6800 0.7725 ;
        RECT 1.0500 0.2775 1.1775 0.3975 ;
        RECT 1.0500 0.6525 1.1775 0.7725 ;
    END
END CKN_0101


MACRO CKN_0110
    CLASS CORE ;
    FOREIGN CKN_0110 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.4700 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 0.8925 0.2775 1.0500 0.3975 ;
        RECT 0.8925 0.6525 1.0500 0.7725 ;
        RECT 0.5775 0.2775 0.8925 0.7725 ;
        RECT 0.4200 0.2775 0.5775 0.3975 ;
        RECT 0.4200 0.6525 0.5775 0.7725 ;
        VIA 0.8925 0.3375 VIA12_slot ;
        VIA 0.8925 0.7125 VIA12_slot ;
        VIA 0.5775 0.3375 VIA12_slot ;
        VIA 0.5775 0.7125 VIA12_slot ;
        END
    END ZN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1425 0.4725 1.3350 0.5475 ;
        RECT 0.0675 0.3675 0.1425 0.6825 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.4250 -0.0750 1.4700 0.0750 ;
        RECT 1.3050 -0.0750 1.4250 0.2925 ;
        RECT 1.0050 -0.0750 1.3050 0.0750 ;
        RECT 0.8850 -0.0750 1.0050 0.2025 ;
        RECT 0.5850 -0.0750 0.8850 0.0750 ;
        RECT 0.4650 -0.0750 0.5850 0.2025 ;
        RECT 0.1425 -0.0750 0.4650 0.0750 ;
        RECT 0.0675 -0.0750 0.1425 0.2475 ;
        RECT 0.0000 -0.0750 0.0675 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.4250 0.9750 1.4700 1.1250 ;
        RECT 1.3050 0.6600 1.4250 1.1250 ;
        RECT 1.0050 0.9750 1.3050 1.1250 ;
        RECT 0.8850 0.8475 1.0050 1.1250 ;
        RECT 0.5850 0.9750 0.8850 1.1250 ;
        RECT 0.4650 0.8475 0.5850 1.1250 ;
        RECT 0.1425 0.9750 0.4650 1.1250 ;
        RECT 0.0675 0.8025 0.1425 1.1250 ;
        RECT 0.0000 0.9750 0.0675 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.3350 0.2250 1.3950 0.2850 ;
        RECT 1.3350 0.6675 1.3950 0.7275 ;
        RECT 1.3350 0.8325 1.3950 0.8925 ;
        RECT 1.2300 0.4800 1.2900 0.5400 ;
        RECT 1.1250 0.2700 1.1850 0.3300 ;
        RECT 1.1250 0.6825 1.1850 0.7425 ;
        RECT 1.0200 0.4800 1.0800 0.5400 ;
        RECT 0.9150 0.1350 0.9750 0.1950 ;
        RECT 0.9150 0.8550 0.9750 0.9150 ;
        RECT 0.8100 0.4800 0.8700 0.5400 ;
        RECT 0.7050 0.2700 0.7650 0.3300 ;
        RECT 0.7050 0.6825 0.7650 0.7425 ;
        RECT 0.6000 0.4800 0.6600 0.5400 ;
        RECT 0.4950 0.1350 0.5550 0.1950 ;
        RECT 0.4950 0.8550 0.5550 0.9150 ;
        RECT 0.3900 0.4800 0.4500 0.5400 ;
        RECT 0.2850 0.2700 0.3450 0.3300 ;
        RECT 0.2850 0.6825 0.3450 0.7425 ;
        RECT 0.1800 0.4800 0.2400 0.5400 ;
        RECT 0.0750 0.1575 0.1350 0.2175 ;
        RECT 0.0750 0.8325 0.1350 0.8925 ;
        LAYER M1 ;
        RECT 1.0950 0.2400 1.2150 0.3975 ;
        RECT 0.2775 0.6525 1.2000 0.7725 ;
        RECT 0.7950 0.2775 1.0950 0.3975 ;
        RECT 0.6750 0.2400 0.7950 0.3975 ;
        RECT 0.3750 0.2775 0.6750 0.3975 ;
        RECT 0.2550 0.2400 0.3750 0.3975 ;
        LAYER M2 ;
        RECT 0.9225 0.2775 1.0500 0.3975 ;
        RECT 0.9225 0.6525 1.0500 0.7725 ;
        RECT 0.4200 0.2775 0.5475 0.3975 ;
        RECT 0.4200 0.6525 0.5475 0.7725 ;
    END
END CKN_0110


MACRO CKN_0111
    CLASS CORE ;
    FOREIGN CKN_0111 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.0500 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 0.3675 0.2700 0.6825 0.7800 ;
        VIA 0.5250 0.3525 VIA12_slot ;
        VIA 0.5250 0.6975 VIA12_slot ;
        END
    END ZN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1425 0.4725 0.9150 0.5475 ;
        RECT 0.0675 0.3675 0.1425 0.6825 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.0050 -0.0750 1.0500 0.0750 ;
        RECT 0.8850 -0.0750 1.0050 0.2925 ;
        RECT 0.5850 -0.0750 0.8850 0.0750 ;
        RECT 0.4650 -0.0750 0.5850 0.2025 ;
        RECT 0.1425 -0.0750 0.4650 0.0750 ;
        RECT 0.0675 -0.0750 0.1425 0.2475 ;
        RECT 0.0000 -0.0750 0.0675 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.0050 0.9750 1.0500 1.1250 ;
        RECT 0.8850 0.6600 1.0050 1.1250 ;
        RECT 0.5850 0.9750 0.8850 1.1250 ;
        RECT 0.4650 0.8475 0.5850 1.1250 ;
        RECT 0.1425 0.9750 0.4650 1.1250 ;
        RECT 0.0675 0.8025 0.1425 1.1250 ;
        RECT 0.0000 0.9750 0.0675 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 0.9150 0.2175 0.9750 0.2775 ;
        RECT 0.9150 0.6675 0.9750 0.7275 ;
        RECT 0.9150 0.8325 0.9750 0.8925 ;
        RECT 0.8100 0.4800 0.8700 0.5400 ;
        RECT 0.7050 0.2325 0.7650 0.2925 ;
        RECT 0.7050 0.6825 0.7650 0.7425 ;
        RECT 0.6000 0.4800 0.6600 0.5400 ;
        RECT 0.4950 0.1350 0.5550 0.1950 ;
        RECT 0.4950 0.8550 0.5550 0.9150 ;
        RECT 0.3900 0.4800 0.4500 0.5400 ;
        RECT 0.2850 0.2325 0.3450 0.2925 ;
        RECT 0.2850 0.6825 0.3450 0.7425 ;
        RECT 0.1800 0.4800 0.2400 0.5400 ;
        RECT 0.0750 0.1575 0.1350 0.2175 ;
        RECT 0.0750 0.8325 0.1350 0.8925 ;
        LAYER M1 ;
        RECT 0.6750 0.2025 0.7950 0.3975 ;
        RECT 0.2775 0.6525 0.7800 0.7725 ;
        RECT 0.3750 0.2775 0.6750 0.3975 ;
        RECT 0.2550 0.2025 0.3750 0.3975 ;
    END
END CKN_0111


MACRO CKN_1000
    CLASS CORE ;
    FOREIGN CKN_1000 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.4200 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.3075 0.1500 0.3825 0.8475 ;
        RECT 0.2550 0.1500 0.3075 0.2550 ;
        RECT 0.2775 0.6675 0.3075 0.8475 ;
        END
    END ZN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1425 0.4425 0.2325 0.5925 ;
        RECT 0.0675 0.3675 0.1425 0.6825 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.1650 -0.0750 0.4200 0.0750 ;
        RECT 0.0450 -0.0750 0.1650 0.2325 ;
        RECT 0.0000 -0.0750 0.0450 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.1650 0.9750 0.4200 1.1250 ;
        RECT 0.0450 0.8100 0.1650 1.1250 ;
        RECT 0.0000 0.9750 0.0450 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 0.2850 0.1575 0.3450 0.2175 ;
        RECT 0.2850 0.7575 0.3450 0.8175 ;
        RECT 0.1725 0.4875 0.2325 0.5475 ;
        RECT 0.0750 0.1575 0.1350 0.2175 ;
        RECT 0.0750 0.8250 0.1350 0.8850 ;
    END
END CKN_1000


MACRO CKN_1010
    CLASS CORE ;
    FOREIGN CKN_1010 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.4200 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.3075 0.2025 0.3825 0.8475 ;
        RECT 0.2775 0.2025 0.3075 0.3825 ;
        RECT 0.2775 0.6675 0.3075 0.8475 ;
        END
    END ZN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1425 0.4425 0.2325 0.5925 ;
        RECT 0.0675 0.3675 0.1425 0.6825 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.1425 -0.0750 0.4200 0.0750 ;
        RECT 0.0675 -0.0750 0.1425 0.2475 ;
        RECT 0.0000 -0.0750 0.0675 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.1425 0.9750 0.4200 1.1250 ;
        RECT 0.0675 0.8025 0.1425 1.1250 ;
        RECT 0.0000 0.9750 0.0675 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 0.2850 0.2325 0.3450 0.2925 ;
        RECT 0.2850 0.7425 0.3450 0.8025 ;
        RECT 0.1725 0.4875 0.2325 0.5475 ;
        RECT 0.0750 0.1575 0.1350 0.2175 ;
        RECT 0.0750 0.8325 0.1350 0.8925 ;
    END
END CKN_1010


MACRO CKN_1100
    CLASS CORE ;
    FOREIGN CKN_1100 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.5700 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 1.9425 0.2775 2.1000 0.3975 ;
        RECT 1.9425 0.6525 2.1000 0.7725 ;
        RECT 1.6275 0.2775 1.9425 0.7725 ;
        RECT 1.4700 0.2775 1.6275 0.3975 ;
        RECT 1.4700 0.6525 1.6275 0.7725 ;
        VIA 1.9425 0.3375 VIA12_slot ;
        VIA 1.9425 0.7125 VIA12_slot ;
        VIA 1.6275 0.3375 VIA12_slot ;
        VIA 1.6275 0.7125 VIA12_slot ;
        END
    END ZN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1425 0.4725 3.4650 0.5475 ;
        RECT 0.0675 0.3675 0.1425 0.6825 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 3.5250 -0.0750 3.5700 0.0750 ;
        RECT 3.4050 -0.0750 3.5250 0.2925 ;
        RECT 3.1050 -0.0750 3.4050 0.0750 ;
        RECT 2.9850 -0.0750 3.1050 0.2025 ;
        RECT 2.6850 -0.0750 2.9850 0.0750 ;
        RECT 2.5650 -0.0750 2.6850 0.2025 ;
        RECT 2.2650 -0.0750 2.5650 0.0750 ;
        RECT 2.1450 -0.0750 2.2650 0.2025 ;
        RECT 1.8450 -0.0750 2.1450 0.0750 ;
        RECT 1.7250 -0.0750 1.8450 0.2025 ;
        RECT 1.4250 -0.0750 1.7250 0.0750 ;
        RECT 1.3050 -0.0750 1.4250 0.2025 ;
        RECT 1.0050 -0.0750 1.3050 0.0750 ;
        RECT 0.8850 -0.0750 1.0050 0.2025 ;
        RECT 0.5850 -0.0750 0.8850 0.0750 ;
        RECT 0.4650 -0.0750 0.5850 0.2025 ;
        RECT 0.1425 -0.0750 0.4650 0.0750 ;
        RECT 0.0675 -0.0750 0.1425 0.2475 ;
        RECT 0.0000 -0.0750 0.0675 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 3.5250 0.9750 3.5700 1.1250 ;
        RECT 3.4050 0.6600 3.5250 1.1250 ;
        RECT 3.1050 0.9750 3.4050 1.1250 ;
        RECT 2.9850 0.8475 3.1050 1.1250 ;
        RECT 2.6850 0.9750 2.9850 1.1250 ;
        RECT 2.5650 0.8475 2.6850 1.1250 ;
        RECT 2.2650 0.9750 2.5650 1.1250 ;
        RECT 2.1450 0.8475 2.2650 1.1250 ;
        RECT 1.8450 0.9750 2.1450 1.1250 ;
        RECT 1.7250 0.8475 1.8450 1.1250 ;
        RECT 1.4250 0.9750 1.7250 1.1250 ;
        RECT 1.3050 0.8475 1.4250 1.1250 ;
        RECT 1.0050 0.9750 1.3050 1.1250 ;
        RECT 0.8850 0.8475 1.0050 1.1250 ;
        RECT 0.5850 0.9750 0.8850 1.1250 ;
        RECT 0.4650 0.8475 0.5850 1.1250 ;
        RECT 0.1425 0.9750 0.4650 1.1250 ;
        RECT 0.0675 0.8025 0.1425 1.1250 ;
        RECT 0.0000 0.9750 0.0675 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 3.4350 0.2250 3.4950 0.2850 ;
        RECT 3.4350 0.6675 3.4950 0.7275 ;
        RECT 3.4350 0.8325 3.4950 0.8925 ;
        RECT 3.3300 0.4800 3.3900 0.5400 ;
        RECT 3.2250 0.3075 3.2850 0.3675 ;
        RECT 3.2250 0.6825 3.2850 0.7425 ;
        RECT 3.1200 0.4800 3.1800 0.5400 ;
        RECT 3.0150 0.1350 3.0750 0.1950 ;
        RECT 3.0150 0.8550 3.0750 0.9150 ;
        RECT 2.9100 0.4800 2.9700 0.5400 ;
        RECT 2.8050 0.3075 2.8650 0.3675 ;
        RECT 2.8050 0.6825 2.8650 0.7425 ;
        RECT 2.7000 0.4800 2.7600 0.5400 ;
        RECT 2.5950 0.1350 2.6550 0.1950 ;
        RECT 2.5950 0.8550 2.6550 0.9150 ;
        RECT 2.4900 0.4800 2.5500 0.5400 ;
        RECT 2.3850 0.3075 2.4450 0.3675 ;
        RECT 2.3850 0.6825 2.4450 0.7425 ;
        RECT 2.2800 0.4800 2.3400 0.5400 ;
        RECT 2.1750 0.1350 2.2350 0.1950 ;
        RECT 2.1750 0.8550 2.2350 0.9150 ;
        RECT 2.0700 0.4800 2.1300 0.5400 ;
        RECT 1.9650 0.3075 2.0250 0.3675 ;
        RECT 1.9650 0.6825 2.0250 0.7425 ;
        RECT 1.8600 0.4800 1.9200 0.5400 ;
        RECT 1.7550 0.1350 1.8150 0.1950 ;
        RECT 1.7550 0.8550 1.8150 0.9150 ;
        RECT 1.6500 0.4800 1.7100 0.5400 ;
        RECT 1.5450 0.3075 1.6050 0.3675 ;
        RECT 1.5450 0.6825 1.6050 0.7425 ;
        RECT 1.4400 0.4800 1.5000 0.5400 ;
        RECT 1.3350 0.1350 1.3950 0.1950 ;
        RECT 1.3350 0.8550 1.3950 0.9150 ;
        RECT 1.2300 0.4800 1.2900 0.5400 ;
        RECT 1.1250 0.3075 1.1850 0.3675 ;
        RECT 1.1250 0.6825 1.1850 0.7425 ;
        RECT 1.0200 0.4800 1.0800 0.5400 ;
        RECT 0.9150 0.1350 0.9750 0.1950 ;
        RECT 0.9150 0.8550 0.9750 0.9150 ;
        RECT 0.8100 0.4800 0.8700 0.5400 ;
        RECT 0.7050 0.3075 0.7650 0.3675 ;
        RECT 0.7050 0.6825 0.7650 0.7425 ;
        RECT 0.6000 0.4800 0.6600 0.5400 ;
        RECT 0.4950 0.1350 0.5550 0.1950 ;
        RECT 0.4950 0.8550 0.5550 0.9150 ;
        RECT 0.3900 0.4800 0.4500 0.5400 ;
        RECT 0.2850 0.3075 0.3450 0.3675 ;
        RECT 0.2850 0.6825 0.3450 0.7425 ;
        RECT 0.1800 0.4800 0.2400 0.5400 ;
        RECT 0.0750 0.1575 0.1350 0.2175 ;
        RECT 0.0750 0.8325 0.1350 0.8925 ;
        LAYER M1 ;
        RECT 0.2775 0.2775 3.3000 0.3975 ;
        RECT 0.2775 0.6525 3.3000 0.7725 ;
        LAYER M2 ;
        RECT 1.9725 0.2775 2.1000 0.3975 ;
        RECT 1.9725 0.6525 2.1000 0.7725 ;
        RECT 1.4700 0.2775 1.5975 0.3975 ;
        RECT 1.4700 0.6525 1.5975 0.7725 ;
    END
END CKN_1100


MACRO CKXOR2_0011
    CLASS CORE ;
    FOREIGN CKXOR2_0011 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.8900 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 1.7775 0.3075 1.8525 0.7500 ;
        RECT 1.6125 0.3075 1.7775 0.3825 ;
        RECT 1.6125 0.6750 1.7775 0.7500 ;
        RECT 1.5375 0.2175 1.6125 0.3825 ;
        RECT 1.5375 0.6750 1.6125 0.8175 ;
        END
    END Z
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.0950 0.4125 1.5300 0.4875 ;
        RECT 1.0200 0.3750 1.0950 0.4875 ;
        VIA 1.2600 0.4500 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.1350 0.4125 0.6000 0.4875 ;
        VIA 0.3150 0.4500 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.8450 -0.0750 1.8900 0.0750 ;
        RECT 1.7250 -0.0750 1.8450 0.2250 ;
        RECT 1.4025 -0.0750 1.7250 0.0750 ;
        RECT 1.2975 -0.0750 1.4025 0.2550 ;
        RECT 0.3600 -0.0750 1.2975 0.0750 ;
        RECT 0.2700 -0.0750 0.3600 0.2250 ;
        RECT 0.0000 -0.0750 0.2700 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.8450 0.9750 1.8900 1.1250 ;
        RECT 1.7250 0.8250 1.8450 1.1250 ;
        RECT 1.4250 0.9750 1.7250 1.1250 ;
        RECT 1.3050 0.8700 1.4250 1.1250 ;
        RECT 0.3750 0.9750 1.3050 1.1250 ;
        RECT 0.2550 0.8175 0.3750 1.1250 ;
        RECT 0.0000 0.9750 0.2550 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.7550 0.1575 1.8150 0.2175 ;
        RECT 1.7550 0.8325 1.8150 0.8925 ;
        RECT 1.6425 0.4950 1.7025 0.5550 ;
        RECT 1.5450 0.2925 1.6050 0.3525 ;
        RECT 1.5450 0.7200 1.6050 0.7800 ;
        RECT 1.4400 0.4950 1.5000 0.5550 ;
        RECT 1.3350 0.1650 1.3950 0.2250 ;
        RECT 1.3350 0.8700 1.3950 0.9300 ;
        RECT 1.2300 0.4650 1.2900 0.5250 ;
        RECT 1.1250 0.1575 1.1850 0.2175 ;
        RECT 1.1250 0.7875 1.1850 0.8475 ;
        RECT 1.0125 0.4650 1.0725 0.5250 ;
        RECT 0.9150 0.1575 0.9750 0.2175 ;
        RECT 0.9150 0.8325 0.9750 0.8925 ;
        RECT 0.8100 0.5025 0.8700 0.5625 ;
        RECT 0.7050 0.1800 0.7650 0.2400 ;
        RECT 0.7050 0.8325 0.7650 0.8925 ;
        RECT 0.6075 0.6300 0.6675 0.6900 ;
        RECT 0.3900 0.3450 0.4500 0.4050 ;
        RECT 0.3900 0.6225 0.4500 0.6825 ;
        RECT 0.2850 0.1350 0.3450 0.1950 ;
        RECT 0.2850 0.8400 0.3450 0.9000 ;
        RECT 0.1875 0.4425 0.2475 0.5025 ;
        RECT 0.0750 0.1800 0.1350 0.2400 ;
        RECT 0.0750 0.8325 0.1350 0.8925 ;
        LAYER M1 ;
        RECT 1.4625 0.4650 1.7025 0.5850 ;
        RECT 1.3725 0.4650 1.4625 0.7950 ;
        RECT 1.3050 0.6300 1.3725 0.7950 ;
        RECT 1.1475 0.3300 1.2975 0.5550 ;
        RECT 0.8775 0.1500 1.2225 0.2550 ;
        RECT 1.1100 0.6600 1.2150 0.8850 ;
        RECT 0.6975 0.6600 1.1100 0.7350 ;
        RECT 0.9975 0.3300 1.0725 0.5550 ;
        RECT 0.6300 0.8100 1.0050 0.9000 ;
        RECT 0.3525 0.3300 0.9975 0.4050 ;
        RECT 0.7725 0.4800 0.8925 0.5850 ;
        RECT 0.4950 0.1500 0.7950 0.2550 ;
        RECT 0.5025 0.4800 0.7725 0.5550 ;
        RECT 0.5775 0.6300 0.6975 0.7350 ;
        RECT 0.4275 0.4800 0.5025 0.6975 ;
        RECT 0.1650 0.6225 0.4275 0.6975 ;
        RECT 0.2775 0.3300 0.3525 0.5325 ;
        RECT 0.1875 0.4125 0.2775 0.5325 ;
        RECT 0.1125 0.6225 0.1650 0.9000 ;
        RECT 0.1125 0.1500 0.1425 0.2700 ;
        RECT 0.0375 0.1500 0.1125 0.9000 ;
        LAYER VIA1 ;
        RECT 1.3050 0.6750 1.3800 0.7500 ;
        RECT 0.9450 0.6600 1.0200 0.7350 ;
        RECT 0.9225 0.1650 0.9975 0.2400 ;
        RECT 0.7650 0.8100 0.8400 0.8850 ;
        RECT 0.6825 0.1650 0.7575 0.2400 ;
        LAYER M2 ;
        RECT 1.2900 0.6300 1.3950 0.8850 ;
        RECT 0.7950 0.8100 1.2900 0.8850 ;
        RECT 0.9450 0.6600 1.0650 0.7350 ;
        RECT 0.9450 0.1500 1.0425 0.2550 ;
        RECT 0.8700 0.1500 0.9450 0.7350 ;
        RECT 0.7200 0.1500 0.7950 0.8850 ;
        RECT 0.6450 0.1500 0.7200 0.2550 ;
    END
END CKXOR2_0011


MACRO CKXOR2_0111
    CLASS CORE ;
    FOREIGN CKXOR2_0111 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.3600 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 2.6775 0.2400 2.9925 0.7500 ;
        VIA 2.8350 0.3225 VIA12_slot ;
        VIA 2.8350 0.6675 VIA12_slot ;
        END
    END Z
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 2.0775 0.4425 2.1525 0.6375 ;
        RECT 1.6125 0.5625 2.0775 0.6375 ;
        VIA 2.1150 0.5250 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.6275 0.4125 1.7775 0.4875 ;
        RECT 1.5525 0.3225 1.6275 0.4875 ;
        RECT 1.0950 0.3225 1.5525 0.4050 ;
        RECT 1.0200 0.3225 1.0950 0.4875 ;
        RECT 0.4725 0.4125 1.0200 0.4875 ;
        RECT 0.3675 0.2625 0.4725 0.4875 ;
        VIA 1.6650 0.4500 VIA12_square ;
        VIA 0.9525 0.4500 VIA12_square ;
        VIA 0.4200 0.3375 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 3.2925 -0.0750 3.3600 0.0750 ;
        RECT 3.2175 -0.0750 3.2925 0.3150 ;
        RECT 2.8950 -0.0750 3.2175 0.0750 ;
        RECT 2.7750 -0.0750 2.8950 0.1950 ;
        RECT 2.4525 -0.0750 2.7750 0.0750 ;
        RECT 2.3775 -0.0750 2.4525 0.3075 ;
        RECT 2.0625 -0.0750 2.3775 0.0750 ;
        RECT 1.9575 -0.0750 2.0625 0.2475 ;
        RECT 1.0050 -0.0750 1.9575 0.0750 ;
        RECT 0.8850 -0.0750 1.0050 0.1875 ;
        RECT 0.3750 -0.0750 0.8850 0.0750 ;
        RECT 0.2550 -0.0750 0.3750 0.2250 ;
        RECT 0.0000 -0.0750 0.2550 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 3.2925 0.9750 3.3600 1.1250 ;
        RECT 3.2175 0.7200 3.2925 1.1250 ;
        RECT 2.8875 0.9750 3.2175 1.1250 ;
        RECT 2.7825 0.8025 2.8875 1.1250 ;
        RECT 2.4750 0.9750 2.7825 1.1250 ;
        RECT 2.3550 0.8025 2.4750 1.1250 ;
        RECT 2.0550 0.9750 2.3550 1.1250 ;
        RECT 1.9350 0.8025 2.0550 1.1250 ;
        RECT 0.7875 0.9750 1.9350 1.1250 ;
        RECT 0.6825 0.7875 0.7875 1.1250 ;
        RECT 0.3675 0.9750 0.6825 1.1250 ;
        RECT 0.2625 0.8100 0.3675 1.1250 ;
        RECT 0.0000 0.9750 0.2625 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 3.2250 0.2250 3.2850 0.2850 ;
        RECT 3.2250 0.7650 3.2850 0.8250 ;
        RECT 3.1200 0.4650 3.1800 0.5250 ;
        RECT 3.0150 0.2250 3.0750 0.2850 ;
        RECT 3.0150 0.7575 3.0750 0.8175 ;
        RECT 2.9100 0.4650 2.9700 0.5250 ;
        RECT 2.8050 0.1275 2.8650 0.1875 ;
        RECT 2.8050 0.8325 2.8650 0.8925 ;
        RECT 2.7000 0.4650 2.7600 0.5250 ;
        RECT 2.5950 0.2250 2.6550 0.2850 ;
        RECT 2.5950 0.7575 2.6550 0.8175 ;
        RECT 2.4900 0.4650 2.5500 0.5250 ;
        RECT 2.3850 0.2175 2.4450 0.2775 ;
        RECT 2.3850 0.8325 2.4450 0.8925 ;
        RECT 2.2800 0.4875 2.3400 0.5475 ;
        RECT 2.1750 0.1950 2.2350 0.2550 ;
        RECT 2.1750 0.7725 2.2350 0.8325 ;
        RECT 2.0700 0.4875 2.1300 0.5475 ;
        RECT 1.9650 0.1575 2.0250 0.2175 ;
        RECT 1.9650 0.8100 2.0250 0.8700 ;
        RECT 1.7550 0.7725 1.8150 0.8325 ;
        RECT 1.6500 0.4500 1.7100 0.5100 ;
        RECT 1.5450 0.1725 1.6050 0.2325 ;
        RECT 1.5450 0.8250 1.6050 0.8850 ;
        RECT 1.4400 0.4725 1.5000 0.5325 ;
        RECT 1.3350 0.2175 1.3950 0.2775 ;
        RECT 1.3350 0.8175 1.3950 0.8775 ;
        RECT 1.2300 0.6300 1.2900 0.6900 ;
        RECT 1.1250 0.2100 1.1850 0.2700 ;
        RECT 1.1250 0.8175 1.1850 0.8775 ;
        RECT 1.0200 0.4650 1.0800 0.5250 ;
        RECT 0.9150 0.1275 0.9750 0.1875 ;
        RECT 0.8100 0.4650 0.8700 0.5250 ;
        RECT 0.7050 0.1875 0.7650 0.2475 ;
        RECT 0.7050 0.8175 0.7650 0.8775 ;
        RECT 0.6000 0.4800 0.6600 0.5400 ;
        RECT 0.4950 0.8175 0.5550 0.8775 ;
        RECT 0.3900 0.4800 0.4500 0.5400 ;
        RECT 0.2850 0.1575 0.3450 0.2175 ;
        RECT 0.2850 0.8325 0.3450 0.8925 ;
        RECT 0.1875 0.4725 0.2475 0.5325 ;
        RECT 0.0750 0.1650 0.1350 0.2250 ;
        RECT 0.0750 0.8325 0.1350 0.8925 ;
        LAYER M1 ;
        RECT 2.4375 0.4425 3.2100 0.5475 ;
        RECT 2.9925 0.1950 3.0975 0.3675 ;
        RECT 3.0075 0.6225 3.0825 0.8700 ;
        RECT 2.6625 0.6225 3.0075 0.7125 ;
        RECT 2.6775 0.2775 2.9925 0.3675 ;
        RECT 2.5725 0.1950 2.6775 0.3675 ;
        RECT 2.5875 0.6225 2.6625 0.8700 ;
        RECT 2.2575 0.4650 2.3625 0.5700 ;
        RECT 2.1900 0.1725 2.2650 0.3900 ;
        RECT 1.9950 0.4800 2.2575 0.5700 ;
        RECT 2.1675 0.6450 2.2425 0.8700 ;
        RECT 2.1450 0.1725 2.1900 0.3975 ;
        RECT 1.8825 0.6450 2.1675 0.7200 ;
        RECT 1.8825 0.3225 2.1450 0.3975 ;
        RECT 1.8225 0.1500 1.8825 0.7200 ;
        RECT 1.8075 0.1500 1.8225 0.8625 ;
        RECT 1.5225 0.1500 1.8075 0.2550 ;
        RECT 1.7475 0.6450 1.8075 0.8625 ;
        RECT 1.4850 0.6450 1.7475 0.7200 ;
        RECT 1.5975 0.3300 1.7325 0.5700 ;
        RECT 1.3125 0.7950 1.6575 0.9000 ;
        RECT 1.2075 0.4500 1.5225 0.5550 ;
        RECT 1.4250 0.6300 1.4850 0.7200 ;
        RECT 1.2675 0.1500 1.4250 0.3600 ;
        RECT 1.1925 0.6300 1.4250 0.7050 ;
        RECT 1.0875 0.7950 1.2075 0.9000 ;
        RECT 1.1175 0.1800 1.1925 0.3375 ;
        RECT 0.7950 0.2625 1.1175 0.3375 ;
        RECT 1.0125 0.6375 1.0875 0.9000 ;
        RECT 0.8100 0.4125 1.0800 0.5550 ;
        RECT 0.6075 0.6375 1.0125 0.7125 ;
        RECT 0.6750 0.1800 0.7950 0.3375 ;
        RECT 0.4575 0.4500 0.6900 0.5550 ;
        RECT 0.5325 0.6375 0.6075 0.9000 ;
        RECT 0.4725 0.7950 0.5325 0.9000 ;
        RECT 0.3075 0.3000 0.5025 0.3750 ;
        RECT 0.3825 0.4500 0.4575 0.7200 ;
        RECT 0.1650 0.6450 0.3825 0.7200 ;
        RECT 0.2325 0.3000 0.3075 0.5625 ;
        RECT 0.1875 0.4425 0.2325 0.5625 ;
        RECT 0.1125 0.1500 0.1650 0.2625 ;
        RECT 0.1125 0.6450 0.1650 0.9000 ;
        RECT 0.0375 0.1500 0.1125 0.9000 ;
        LAYER VIA1 ;
        RECT 2.4750 0.4575 2.5500 0.5325 ;
        RECT 1.4625 0.8100 1.5375 0.8850 ;
        RECT 1.3125 0.1650 1.3875 0.2400 ;
        RECT 1.2750 0.4800 1.3500 0.5550 ;
        RECT 0.3825 0.5625 0.4575 0.6375 ;
        LAYER M2 ;
        RECT 2.3325 0.4200 2.5650 0.5700 ;
        RECT 2.2575 0.1650 2.3325 0.8850 ;
        RECT 1.2675 0.1650 2.2575 0.2400 ;
        RECT 1.4175 0.8100 2.2575 0.8850 ;
        RECT 1.2600 0.4800 1.4025 0.5550 ;
        RECT 1.1850 0.4800 1.2600 0.6375 ;
        RECT 0.3075 0.5625 1.1850 0.6375 ;
    END
END CKXOR2_0111


MACRO CKXOR2_1000
    CLASS CORE ;
    FOREIGN CKXOR2_1000 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.6800 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 1.5675 0.1500 1.6425 0.9000 ;
        RECT 1.5150 0.1500 1.5675 0.3825 ;
        RECT 1.5225 0.6675 1.5675 0.9000 ;
        RECT 1.5000 0.7950 1.5225 0.9000 ;
        END
    END Z
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.1475 0.1125 1.6200 0.1875 ;
        RECT 1.1475 0.4125 1.2750 0.4875 ;
        RECT 1.0725 0.1125 1.1475 0.4875 ;
        VIA 1.1925 0.4500 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.1200 0.4125 0.5850 0.4875 ;
        VIA 0.2925 0.4500 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.4025 -0.0750 1.6800 0.0750 ;
        RECT 1.2975 -0.0750 1.4025 0.2475 ;
        RECT 0.3750 -0.0750 1.2975 0.0750 ;
        RECT 0.2550 -0.0750 0.3750 0.2250 ;
        RECT 0.0000 -0.0750 0.2550 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.4250 0.9750 1.6800 1.1250 ;
        RECT 1.3050 0.8325 1.4250 1.1250 ;
        RECT 0.3750 0.9750 1.3050 1.1250 ;
        RECT 0.2550 0.8325 0.3750 1.1250 ;
        RECT 0.0000 0.9750 0.2550 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.5450 0.1575 1.6050 0.2175 ;
        RECT 1.5450 0.8325 1.6050 0.8925 ;
        RECT 1.4325 0.4875 1.4925 0.5475 ;
        RECT 1.3350 0.1575 1.3950 0.2175 ;
        RECT 1.3350 0.8325 1.3950 0.8925 ;
        RECT 1.2300 0.4650 1.2900 0.5250 ;
        RECT 1.1250 0.1575 1.1850 0.2175 ;
        RECT 1.1250 0.8100 1.1850 0.8700 ;
        RECT 1.0125 0.4650 1.0725 0.5250 ;
        RECT 0.9150 0.1575 0.9750 0.2175 ;
        RECT 0.9150 0.8325 0.9750 0.8925 ;
        RECT 0.8100 0.5025 0.8700 0.5625 ;
        RECT 0.7050 0.1800 0.7650 0.2400 ;
        RECT 0.7050 0.8325 0.7650 0.8925 ;
        RECT 0.6000 0.6525 0.6600 0.7125 ;
        RECT 0.3975 0.6600 0.4575 0.7200 ;
        RECT 0.3900 0.3450 0.4500 0.4050 ;
        RECT 0.2850 0.1575 0.3450 0.2175 ;
        RECT 0.2850 0.8325 0.3450 0.8925 ;
        RECT 0.1875 0.4800 0.2475 0.5400 ;
        RECT 0.0750 0.1575 0.1350 0.2175 ;
        RECT 0.0750 0.8175 0.1350 0.8775 ;
        LAYER M1 ;
        RECT 1.4475 0.4575 1.4925 0.5775 ;
        RECT 1.3725 0.4575 1.4475 0.7350 ;
        RECT 1.2900 0.6300 1.3725 0.7350 ;
        RECT 1.1475 0.3300 1.2975 0.5550 ;
        RECT 0.8700 0.1500 1.2225 0.2550 ;
        RECT 1.1100 0.6600 1.2150 0.9000 ;
        RECT 0.6825 0.6600 1.1100 0.7350 ;
        RECT 0.9975 0.3300 1.0725 0.5550 ;
        RECT 0.5775 0.8100 1.0050 0.9000 ;
        RECT 0.3450 0.3300 0.9975 0.4050 ;
        RECT 0.7725 0.4800 0.8925 0.5850 ;
        RECT 0.4725 0.1500 0.7950 0.2550 ;
        RECT 0.5025 0.4800 0.7725 0.5550 ;
        RECT 0.5775 0.6300 0.6825 0.7350 ;
        RECT 0.4275 0.4800 0.5025 0.7275 ;
        RECT 0.1575 0.6525 0.4275 0.7275 ;
        RECT 0.2325 0.3300 0.3450 0.5775 ;
        RECT 0.1875 0.4500 0.2325 0.5775 ;
        RECT 0.1125 0.1500 0.1650 0.2700 ;
        RECT 0.1125 0.6525 0.1575 0.9000 ;
        RECT 0.0375 0.1500 0.1125 0.9000 ;
        LAYER VIA1 ;
        RECT 1.3725 0.5625 1.4475 0.6375 ;
        RECT 0.9375 0.6600 1.0125 0.7350 ;
        RECT 0.9075 0.1650 0.9825 0.2400 ;
        RECT 0.7500 0.8100 0.8250 0.8850 ;
        RECT 0.6675 0.1650 0.7425 0.2400 ;
        LAYER M2 ;
        RECT 1.2900 0.5625 1.5225 0.6375 ;
        RECT 1.2150 0.5625 1.2900 0.8850 ;
        RECT 0.7800 0.8100 1.2150 0.8850 ;
        RECT 0.9675 0.6600 1.0575 0.7350 ;
        RECT 0.9675 0.1275 0.9975 0.2775 ;
        RECT 0.8925 0.1275 0.9675 0.7350 ;
        RECT 0.7050 0.1500 0.7800 0.8850 ;
        RECT 0.6300 0.1500 0.7050 0.2550 ;
    END
END CKXOR2_1000


MACRO CKXOR2_1010
    CLASS CORE ;
    FOREIGN CKXOR2_1010 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.6800 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 1.5675 0.2175 1.6425 0.8325 ;
        RECT 1.5375 0.2175 1.5675 0.3825 ;
        RECT 1.5375 0.6675 1.5675 0.8325 ;
        END
    END Z
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.0950 0.4125 1.5450 0.4875 ;
        RECT 1.0200 0.3750 1.0950 0.4875 ;
        VIA 1.2600 0.4500 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.1350 0.4125 0.6000 0.4875 ;
        VIA 0.3150 0.4500 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.4250 -0.0750 1.6800 0.0750 ;
        RECT 1.3050 -0.0750 1.4250 0.2175 ;
        RECT 0.3750 -0.0750 1.3050 0.0750 ;
        RECT 0.2550 -0.0750 0.3750 0.2250 ;
        RECT 0.0000 -0.0750 0.2550 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.4250 0.9750 1.6800 1.1250 ;
        RECT 1.3200 0.8400 1.4250 1.1250 ;
        RECT 0.3750 0.9750 1.3200 1.1250 ;
        RECT 0.2550 0.8175 0.3750 1.1250 ;
        RECT 0.0000 0.9750 0.2550 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.5450 0.2700 1.6050 0.3300 ;
        RECT 1.5450 0.7350 1.6050 0.7950 ;
        RECT 1.4325 0.4950 1.4925 0.5550 ;
        RECT 1.3350 0.1275 1.3950 0.1875 ;
        RECT 1.3350 0.8700 1.3950 0.9300 ;
        RECT 1.2225 0.4500 1.2825 0.5100 ;
        RECT 1.1250 0.1575 1.1850 0.2175 ;
        RECT 1.1250 0.8325 1.1850 0.8925 ;
        RECT 1.0200 0.4500 1.0800 0.5100 ;
        RECT 0.9150 0.1575 0.9750 0.2175 ;
        RECT 0.9150 0.8325 0.9750 0.8925 ;
        RECT 0.8025 0.4875 0.8625 0.5475 ;
        RECT 0.7050 0.1800 0.7650 0.2400 ;
        RECT 0.7050 0.8325 0.7650 0.8925 ;
        RECT 0.6000 0.6525 0.6600 0.7125 ;
        RECT 0.3900 0.3450 0.4500 0.4050 ;
        RECT 0.3900 0.6525 0.4500 0.7125 ;
        RECT 0.2850 0.1350 0.3450 0.1950 ;
        RECT 0.2850 0.8400 0.3450 0.9000 ;
        RECT 0.1875 0.4800 0.2475 0.5400 ;
        RECT 0.0750 0.1800 0.1350 0.2400 ;
        RECT 0.0750 0.8175 0.1350 0.8775 ;
        LAYER M1 ;
        RECT 1.4625 0.4650 1.4925 0.5850 ;
        RECT 1.3875 0.4650 1.4625 0.7500 ;
        RECT 1.3125 0.3150 1.4325 0.3900 ;
        RECT 1.2375 0.6000 1.3875 0.7500 ;
        RECT 1.2675 0.3150 1.3125 0.5250 ;
        RECT 1.1775 0.3300 1.2675 0.5250 ;
        RECT 0.8775 0.1500 1.2150 0.2550 ;
        RECT 1.1550 0.8250 1.2150 0.9000 ;
        RECT 1.0800 0.6300 1.1550 0.9000 ;
        RECT 0.9975 0.3300 1.1025 0.5400 ;
        RECT 0.6900 0.6300 1.0800 0.7050 ;
        RECT 0.8625 0.7950 1.0050 0.9000 ;
        RECT 0.3525 0.3300 0.9975 0.4050 ;
        RECT 0.5025 0.4800 0.8925 0.5550 ;
        RECT 0.6300 0.8100 0.8625 0.9000 ;
        RECT 0.4950 0.1500 0.7950 0.2550 ;
        RECT 0.5775 0.6300 0.6900 0.7350 ;
        RECT 0.4275 0.4800 0.5025 0.7200 ;
        RECT 0.1575 0.6450 0.4275 0.7200 ;
        RECT 0.2775 0.3300 0.3525 0.5700 ;
        RECT 0.1875 0.4500 0.2775 0.5700 ;
        RECT 0.1125 0.6450 0.1575 0.9000 ;
        RECT 0.1125 0.1500 0.1425 0.2700 ;
        RECT 0.0375 0.1500 0.1125 0.9000 ;
        LAYER VIA1 ;
        RECT 1.2525 0.6375 1.3275 0.7125 ;
        RECT 0.9300 0.6300 1.0050 0.7050 ;
        RECT 0.9225 0.1650 0.9975 0.2400 ;
        RECT 0.7650 0.8100 0.8400 0.8850 ;
        RECT 0.6825 0.1650 0.7575 0.2400 ;
        LAYER M2 ;
        RECT 1.2225 0.5775 1.3275 0.8850 ;
        RECT 0.7950 0.8100 1.2225 0.8850 ;
        RECT 0.9450 0.6300 1.0800 0.7050 ;
        RECT 0.9450 0.1500 1.0425 0.2550 ;
        RECT 0.8700 0.1500 0.9450 0.7050 ;
        RECT 0.7200 0.1500 0.7950 0.8850 ;
        RECT 0.6450 0.1500 0.7200 0.2550 ;
    END
END CKXOR2_1010


MACRO DCAP16_0010
    CLASS CORE ;
    FOREIGN DCAP16_0010 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.3600 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.1575 -0.0750 3.3600 0.0750 ;
        RECT 0.0525 -0.0750 0.1575 0.2625 ;
        RECT 0.0000 -0.0750 0.0525 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 3.3075 0.9750 3.3600 1.1250 ;
        RECT 3.2025 0.7725 3.3075 1.1250 ;
        RECT 3.0975 0.9750 3.2025 1.1250 ;
        RECT 2.9925 0.7725 3.0975 1.1250 ;
        RECT 2.8875 0.9750 2.9925 1.1250 ;
        RECT 2.7825 0.7725 2.8875 1.1250 ;
        RECT 2.6775 0.9750 2.7825 1.1250 ;
        RECT 2.5725 0.7725 2.6775 1.1250 ;
        RECT 2.4675 0.9750 2.5725 1.1250 ;
        RECT 2.3625 0.7725 2.4675 1.1250 ;
        RECT 2.2575 0.9750 2.3625 1.1250 ;
        RECT 2.1525 0.7725 2.2575 1.1250 ;
        RECT 2.0475 0.9750 2.1525 1.1250 ;
        RECT 1.9425 0.7725 2.0475 1.1250 ;
        RECT 1.8375 0.9750 1.9425 1.1250 ;
        RECT 1.7325 0.7725 1.8375 1.1250 ;
        RECT 1.6275 0.9750 1.7325 1.1250 ;
        RECT 1.5225 0.7725 1.6275 1.1250 ;
        RECT 1.4175 0.9750 1.5225 1.1250 ;
        RECT 1.3125 0.7725 1.4175 1.1250 ;
        RECT 1.2075 0.9750 1.3125 1.1250 ;
        RECT 1.1025 0.7725 1.2075 1.1250 ;
        RECT 0.9975 0.9750 1.1025 1.1250 ;
        RECT 0.8925 0.7725 0.9975 1.1250 ;
        RECT 0.7875 0.9750 0.8925 1.1250 ;
        RECT 0.6825 0.7725 0.7875 1.1250 ;
        RECT 0.5625 0.9750 0.6825 1.1250 ;
        RECT 0.4875 0.7725 0.5625 1.1250 ;
        RECT 0.1575 0.9750 0.4875 1.1250 ;
        RECT 0.0525 0.7725 0.1575 1.1250 ;
        RECT 0.0000 0.9750 0.0525 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 3.2250 0.8025 3.2850 0.8625 ;
        RECT 3.1200 0.6000 3.1800 0.6600 ;
        RECT 3.0150 0.8025 3.0750 0.8625 ;
        RECT 2.9100 0.5475 2.9700 0.6075 ;
        RECT 2.8050 0.8025 2.8650 0.8625 ;
        RECT 2.7000 0.5550 2.7600 0.6150 ;
        RECT 2.5950 0.8025 2.6550 0.8625 ;
        RECT 2.4900 0.5550 2.5500 0.6150 ;
        RECT 2.3850 0.8025 2.4450 0.8625 ;
        RECT 2.2800 0.5550 2.3400 0.6150 ;
        RECT 2.1750 0.8025 2.2350 0.8625 ;
        RECT 2.0700 0.5550 2.1300 0.6150 ;
        RECT 1.9650 0.8025 2.0250 0.8625 ;
        RECT 1.8600 0.5550 1.9200 0.6150 ;
        RECT 1.7550 0.8025 1.8150 0.8625 ;
        RECT 1.6500 0.5550 1.7100 0.6150 ;
        RECT 1.5450 0.8025 1.6050 0.8625 ;
        RECT 1.4400 0.5550 1.5000 0.6150 ;
        RECT 1.3350 0.8025 1.3950 0.8625 ;
        RECT 1.2300 0.5550 1.2900 0.6150 ;
        RECT 1.1250 0.8025 1.1850 0.8625 ;
        RECT 1.0200 0.5550 1.0800 0.6150 ;
        RECT 0.9150 0.8025 0.9750 0.8625 ;
        RECT 0.8100 0.5550 0.8700 0.6150 ;
        RECT 0.7050 0.8025 0.7650 0.8625 ;
        RECT 0.6000 0.5550 0.6600 0.6150 ;
        RECT 0.4950 0.8025 0.5550 0.8625 ;
        RECT 0.2850 0.1800 0.3450 0.2400 ;
        RECT 0.2850 0.7950 0.3450 0.8550 ;
        RECT 0.1800 0.3600 0.2400 0.4200 ;
        RECT 0.1800 0.6000 0.2400 0.6600 ;
        RECT 0.0750 0.1725 0.1350 0.2325 ;
        RECT 0.0750 0.8025 0.1350 0.8625 ;
        LAYER M1 ;
        RECT 3.0900 0.5400 3.2100 0.6600 ;
        RECT 0.7125 0.5400 3.0900 0.6150 ;
        RECT 0.6750 0.5400 0.7125 0.6525 ;
        RECT 0.6000 0.1575 0.6750 0.6525 ;
        RECT 0.2625 0.1575 0.6000 0.2625 ;
        RECT 0.5475 0.5400 0.6000 0.6525 ;
        RECT 0.1425 0.3525 0.3375 0.4275 ;
        RECT 0.2550 0.7725 0.3375 0.8775 ;
        RECT 0.0975 0.5025 0.2625 0.6975 ;
        RECT 0.3375 0.3525 0.4125 0.8775 ;
        LAYER VIA1 ;
        RECT 0.5850 0.5625 0.6600 0.6375 ;
        RECT 0.1800 0.5625 0.2550 0.6375 ;
        LAYER M2 ;
        RECT 0.1050 0.5625 0.7350 0.6375 ;
    END
END DCAP16_0010


MACRO DCAP32_0010
    CLASS CORE ;
    FOREIGN DCAP32_0010 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.7200 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.1575 -0.0750 6.7200 0.0750 ;
        RECT 0.0525 -0.0750 0.1575 0.2625 ;
        RECT 0.0000 -0.0750 0.0525 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 6.6675 0.9750 6.7200 1.1250 ;
        RECT 6.5625 0.7725 6.6675 1.1250 ;
        RECT 6.4575 0.9750 6.5625 1.1250 ;
        RECT 6.3525 0.7725 6.4575 1.1250 ;
        RECT 6.2475 0.9750 6.3525 1.1250 ;
        RECT 6.1425 0.7725 6.2475 1.1250 ;
        RECT 6.0375 0.9750 6.1425 1.1250 ;
        RECT 5.9325 0.7725 6.0375 1.1250 ;
        RECT 5.8275 0.9750 5.9325 1.1250 ;
        RECT 5.7225 0.7725 5.8275 1.1250 ;
        RECT 5.6175 0.9750 5.7225 1.1250 ;
        RECT 5.5125 0.7725 5.6175 1.1250 ;
        RECT 5.4075 0.9750 5.5125 1.1250 ;
        RECT 5.3025 0.7725 5.4075 1.1250 ;
        RECT 5.1975 0.9750 5.3025 1.1250 ;
        RECT 5.0925 0.7725 5.1975 1.1250 ;
        RECT 4.9875 0.9750 5.0925 1.1250 ;
        RECT 4.8825 0.7725 4.9875 1.1250 ;
        RECT 4.7775 0.9750 4.8825 1.1250 ;
        RECT 4.6725 0.7725 4.7775 1.1250 ;
        RECT 4.5675 0.9750 4.6725 1.1250 ;
        RECT 4.4625 0.7725 4.5675 1.1250 ;
        RECT 4.3575 0.9750 4.4625 1.1250 ;
        RECT 4.2525 0.7725 4.3575 1.1250 ;
        RECT 4.1475 0.9750 4.2525 1.1250 ;
        RECT 4.0425 0.7725 4.1475 1.1250 ;
        RECT 3.9375 0.9750 4.0425 1.1250 ;
        RECT 3.8325 0.7725 3.9375 1.1250 ;
        RECT 3.7275 0.9750 3.8325 1.1250 ;
        RECT 3.6225 0.7725 3.7275 1.1250 ;
        RECT 3.5175 0.9750 3.6225 1.1250 ;
        RECT 3.4125 0.7725 3.5175 1.1250 ;
        RECT 3.3075 0.9750 3.4125 1.1250 ;
        RECT 3.2025 0.7725 3.3075 1.1250 ;
        RECT 3.0975 0.9750 3.2025 1.1250 ;
        RECT 2.9925 0.7725 3.0975 1.1250 ;
        RECT 2.8875 0.9750 2.9925 1.1250 ;
        RECT 2.7825 0.7725 2.8875 1.1250 ;
        RECT 2.6775 0.9750 2.7825 1.1250 ;
        RECT 2.5725 0.7725 2.6775 1.1250 ;
        RECT 2.4675 0.9750 2.5725 1.1250 ;
        RECT 2.3625 0.7725 2.4675 1.1250 ;
        RECT 2.2575 0.9750 2.3625 1.1250 ;
        RECT 2.1525 0.7725 2.2575 1.1250 ;
        RECT 2.0475 0.9750 2.1525 1.1250 ;
        RECT 1.9425 0.7725 2.0475 1.1250 ;
        RECT 1.8375 0.9750 1.9425 1.1250 ;
        RECT 1.7325 0.7725 1.8375 1.1250 ;
        RECT 1.6275 0.9750 1.7325 1.1250 ;
        RECT 1.5225 0.7725 1.6275 1.1250 ;
        RECT 1.4175 0.9750 1.5225 1.1250 ;
        RECT 1.3125 0.7725 1.4175 1.1250 ;
        RECT 1.2075 0.9750 1.3125 1.1250 ;
        RECT 1.1025 0.7725 1.2075 1.1250 ;
        RECT 0.9975 0.9750 1.1025 1.1250 ;
        RECT 0.8925 0.7725 0.9975 1.1250 ;
        RECT 0.7875 0.9750 0.8925 1.1250 ;
        RECT 0.6825 0.7725 0.7875 1.1250 ;
        RECT 0.5625 0.9750 0.6825 1.1250 ;
        RECT 0.4875 0.7725 0.5625 1.1250 ;
        RECT 0.1575 0.9750 0.4875 1.1250 ;
        RECT 0.0525 0.7725 0.1575 1.1250 ;
        RECT 0.0000 0.9750 0.0525 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 6.5850 0.8025 6.6450 0.8625 ;
        RECT 6.4800 0.6000 6.5400 0.6600 ;
        RECT 6.3750 0.8025 6.4350 0.8625 ;
        RECT 6.2700 0.5475 6.3300 0.6075 ;
        RECT 6.1650 0.8025 6.2250 0.8625 ;
        RECT 6.0600 0.5550 6.1200 0.6150 ;
        RECT 5.9550 0.8025 6.0150 0.8625 ;
        RECT 5.8500 0.5550 5.9100 0.6150 ;
        RECT 5.7450 0.8025 5.8050 0.8625 ;
        RECT 5.6400 0.5550 5.7000 0.6150 ;
        RECT 5.5350 0.8025 5.5950 0.8625 ;
        RECT 5.4300 0.5550 5.4900 0.6150 ;
        RECT 5.3250 0.8025 5.3850 0.8625 ;
        RECT 5.2200 0.5550 5.2800 0.6150 ;
        RECT 5.1150 0.8025 5.1750 0.8625 ;
        RECT 5.0100 0.5550 5.0700 0.6150 ;
        RECT 4.9050 0.8025 4.9650 0.8625 ;
        RECT 4.8000 0.5550 4.8600 0.6150 ;
        RECT 4.6950 0.8025 4.7550 0.8625 ;
        RECT 4.5900 0.5550 4.6500 0.6150 ;
        RECT 4.4850 0.8025 4.5450 0.8625 ;
        RECT 4.3800 0.5550 4.4400 0.6150 ;
        RECT 4.2750 0.8025 4.3350 0.8625 ;
        RECT 4.1700 0.5550 4.2300 0.6150 ;
        RECT 4.0650 0.8025 4.1250 0.8625 ;
        RECT 3.9600 0.5550 4.0200 0.6150 ;
        RECT 3.8550 0.8025 3.9150 0.8625 ;
        RECT 3.7500 0.5550 3.8100 0.6150 ;
        RECT 3.6450 0.8025 3.7050 0.8625 ;
        RECT 3.5400 0.5550 3.6000 0.6150 ;
        RECT 3.4350 0.8025 3.4950 0.8625 ;
        RECT 3.3300 0.5550 3.3900 0.6150 ;
        RECT 3.2250 0.8025 3.2850 0.8625 ;
        RECT 3.1200 0.5550 3.1800 0.6150 ;
        RECT 3.0150 0.8025 3.0750 0.8625 ;
        RECT 2.9100 0.5550 2.9700 0.6150 ;
        RECT 2.8050 0.8025 2.8650 0.8625 ;
        RECT 2.7000 0.5550 2.7600 0.6150 ;
        RECT 2.5950 0.8025 2.6550 0.8625 ;
        RECT 2.4900 0.5550 2.5500 0.6150 ;
        RECT 2.3850 0.8025 2.4450 0.8625 ;
        RECT 0.0750 0.8025 0.1350 0.8625 ;
        RECT 2.2800 0.5550 2.3400 0.6150 ;
        RECT 2.1750 0.8025 2.2350 0.8625 ;
        RECT 2.0700 0.5550 2.1300 0.6150 ;
        RECT 1.9650 0.8025 2.0250 0.8625 ;
        RECT 1.8600 0.5550 1.9200 0.6150 ;
        RECT 1.7550 0.8025 1.8150 0.8625 ;
        RECT 1.6500 0.5550 1.7100 0.6150 ;
        RECT 1.5450 0.8025 1.6050 0.8625 ;
        RECT 1.4400 0.5550 1.5000 0.6150 ;
        RECT 1.3350 0.8025 1.3950 0.8625 ;
        RECT 1.2300 0.5550 1.2900 0.6150 ;
        RECT 1.1250 0.8025 1.1850 0.8625 ;
        RECT 1.0200 0.5550 1.0800 0.6150 ;
        RECT 0.9150 0.8025 0.9750 0.8625 ;
        RECT 0.8100 0.5550 0.8700 0.6150 ;
        RECT 0.7050 0.8025 0.7650 0.8625 ;
        RECT 0.6000 0.5550 0.6600 0.6150 ;
        RECT 0.4950 0.8025 0.5550 0.8625 ;
        RECT 0.2850 0.1800 0.3450 0.2400 ;
        RECT 0.2850 0.8100 0.3450 0.8700 ;
        RECT 0.1800 0.3600 0.2400 0.4200 ;
        RECT 0.1800 0.6000 0.2400 0.6600 ;
        RECT 0.0750 0.1725 0.1350 0.2325 ;
        LAYER M1 ;
        RECT 6.4500 0.5400 6.5700 0.6600 ;
        RECT 0.6825 0.5400 6.4500 0.6150 ;
        RECT 0.6750 0.5400 0.6825 0.6525 ;
        RECT 0.6000 0.1575 0.6750 0.6525 ;
        RECT 0.2625 0.1575 0.6000 0.2625 ;
        RECT 0.5100 0.5400 0.6000 0.6525 ;
        RECT 0.3375 0.3525 0.4125 0.8925 ;
        RECT 0.1425 0.3525 0.3375 0.4275 ;
        RECT 0.2550 0.7875 0.3375 0.8925 ;
        RECT 0.0975 0.5025 0.2625 0.6975 ;
        LAYER VIA1 ;
        RECT 0.5475 0.5625 0.6225 0.6375 ;
        RECT 0.1800 0.5625 0.2550 0.6375 ;
        LAYER M2 ;
        RECT 0.1050 0.5625 0.6975 0.6375 ;
    END
END DCAP32_0010


MACRO DCAP4_0010
    CLASS CORE ;
    FOREIGN DCAP4_0010 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.8400 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.7725 -0.0750 0.8400 0.0750 ;
        RECT 0.6975 -0.0750 0.7725 0.2475 ;
        RECT 0.0000 -0.0750 0.6975 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.7875 0.9750 0.8400 1.1250 ;
        RECT 0.6825 0.7725 0.7875 1.1250 ;
        RECT 0.3525 0.9750 0.6825 1.1250 ;
        RECT 0.2775 0.7725 0.3525 1.1250 ;
        RECT 0.1425 0.9750 0.2775 1.1250 ;
        RECT 0.0675 0.7725 0.1425 1.1250 ;
        RECT 0.0000 0.9750 0.0675 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 0.7050 0.1575 0.7650 0.2175 ;
        RECT 0.7050 0.8025 0.7650 0.8625 ;
        RECT 0.6000 0.3600 0.6600 0.4200 ;
        RECT 0.6000 0.6000 0.6600 0.6600 ;
        RECT 0.4950 0.1875 0.5550 0.2475 ;
        RECT 0.4950 0.7950 0.5550 0.8550 ;
        RECT 0.2850 0.8025 0.3450 0.8625 ;
        RECT 0.1800 0.6000 0.2400 0.6600 ;
        RECT 0.0750 0.8025 0.1350 0.8625 ;
        LAYER M1 ;
        RECT 0.5775 0.5025 0.7650 0.6975 ;
        RECT 0.5025 0.3525 0.7200 0.4275 ;
        RECT 0.1425 0.1800 0.5850 0.2550 ;
        RECT 0.5025 0.7725 0.5850 0.8775 ;
        RECT 0.4275 0.3525 0.5025 0.8775 ;
        RECT 0.1425 0.5325 0.3525 0.6675 ;
        RECT 0.0675 0.1800 0.1425 0.6675 ;
        LAYER VIA1 ;
        RECT 0.5850 0.5625 0.6600 0.6375 ;
        RECT 0.2400 0.5625 0.3150 0.6375 ;
        LAYER M2 ;
        RECT 0.1650 0.5625 0.7350 0.6375 ;
    END
END DCAP4_0010


MACRO DCAP64_0010
    CLASS CORE ;
    FOREIGN DCAP64_0010 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.4400 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 6.6675 -0.0750 13.4400 0.0750 ;
        RECT 6.5625 -0.0750 6.6675 0.2625 ;
        RECT 0.0000 -0.0750 6.5625 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 13.3875 0.9750 13.4400 1.1250 ;
        RECT 13.2825 0.7725 13.3875 1.1250 ;
        RECT 13.1775 0.9750 13.2825 1.1250 ;
        RECT 13.0725 0.7725 13.1775 1.1250 ;
        RECT 12.9675 0.9750 13.0725 1.1250 ;
        RECT 12.8625 0.7725 12.9675 1.1250 ;
        RECT 12.7575 0.9750 12.8625 1.1250 ;
        RECT 12.6525 0.7725 12.7575 1.1250 ;
        RECT 12.5475 0.9750 12.6525 1.1250 ;
        RECT 12.4425 0.7725 12.5475 1.1250 ;
        RECT 12.3375 0.9750 12.4425 1.1250 ;
        RECT 12.2325 0.7725 12.3375 1.1250 ;
        RECT 12.1275 0.9750 12.2325 1.1250 ;
        RECT 12.0225 0.7725 12.1275 1.1250 ;
        RECT 11.9175 0.9750 12.0225 1.1250 ;
        RECT 11.8125 0.7725 11.9175 1.1250 ;
        RECT 11.7075 0.9750 11.8125 1.1250 ;
        RECT 11.6025 0.7725 11.7075 1.1250 ;
        RECT 11.4975 0.9750 11.6025 1.1250 ;
        RECT 11.3925 0.7725 11.4975 1.1250 ;
        RECT 11.2875 0.9750 11.3925 1.1250 ;
        RECT 11.1825 0.7725 11.2875 1.1250 ;
        RECT 11.0775 0.9750 11.1825 1.1250 ;
        RECT 10.9725 0.7725 11.0775 1.1250 ;
        RECT 10.8675 0.9750 10.9725 1.1250 ;
        RECT 10.7625 0.7725 10.8675 1.1250 ;
        RECT 10.6575 0.9750 10.7625 1.1250 ;
        RECT 10.5525 0.7725 10.6575 1.1250 ;
        RECT 10.4475 0.9750 10.5525 1.1250 ;
        RECT 10.3425 0.7725 10.4475 1.1250 ;
        RECT 10.2375 0.9750 10.3425 1.1250 ;
        RECT 10.1325 0.7725 10.2375 1.1250 ;
        RECT 10.0275 0.9750 10.1325 1.1250 ;
        RECT 9.9225 0.7725 10.0275 1.1250 ;
        RECT 9.8175 0.9750 9.9225 1.1250 ;
        RECT 9.7125 0.7725 9.8175 1.1250 ;
        RECT 9.6075 0.9750 9.7125 1.1250 ;
        RECT 9.5025 0.7725 9.6075 1.1250 ;
        RECT 9.3975 0.9750 9.5025 1.1250 ;
        RECT 9.2925 0.7725 9.3975 1.1250 ;
        RECT 9.1875 0.9750 9.2925 1.1250 ;
        RECT 9.0825 0.7725 9.1875 1.1250 ;
        RECT 8.9775 0.9750 9.0825 1.1250 ;
        RECT 8.8725 0.7725 8.9775 1.1250 ;
        RECT 8.7675 0.9750 8.8725 1.1250 ;
        RECT 8.6625 0.7725 8.7675 1.1250 ;
        RECT 8.5575 0.9750 8.6625 1.1250 ;
        RECT 8.4525 0.7725 8.5575 1.1250 ;
        RECT 8.3475 0.9750 8.4525 1.1250 ;
        RECT 8.2425 0.7725 8.3475 1.1250 ;
        RECT 8.1375 0.9750 8.2425 1.1250 ;
        RECT 8.0325 0.7725 8.1375 1.1250 ;
        RECT 7.9275 0.9750 8.0325 1.1250 ;
        RECT 7.8225 0.7725 7.9275 1.1250 ;
        RECT 7.7175 0.9750 7.8225 1.1250 ;
        RECT 7.6125 0.7725 7.7175 1.1250 ;
        RECT 7.5075 0.9750 7.6125 1.1250 ;
        RECT 7.4025 0.7725 7.5075 1.1250 ;
        RECT 7.2975 0.9750 7.4025 1.1250 ;
        RECT 7.1925 0.7725 7.2975 1.1250 ;
        RECT 6.6675 0.9750 7.1925 1.1250 ;
        RECT 6.5625 0.7950 6.6675 1.1250 ;
        RECT 6.4575 0.9750 6.5625 1.1250 ;
        RECT 6.3525 0.7725 6.4575 1.1250 ;
        RECT 6.2475 0.9750 6.3525 1.1250 ;
        RECT 6.1425 0.7725 6.2475 1.1250 ;
        RECT 6.0375 0.9750 6.1425 1.1250 ;
        RECT 5.9325 0.7725 6.0375 1.1250 ;
        RECT 5.8275 0.9750 5.9325 1.1250 ;
        RECT 5.7225 0.7725 5.8275 1.1250 ;
        RECT 5.6175 0.9750 5.7225 1.1250 ;
        RECT 5.5125 0.7725 5.6175 1.1250 ;
        RECT 5.4075 0.9750 5.5125 1.1250 ;
        RECT 5.3025 0.7725 5.4075 1.1250 ;
        RECT 5.1975 0.9750 5.3025 1.1250 ;
        RECT 5.0925 0.7725 5.1975 1.1250 ;
        RECT 4.9875 0.9750 5.0925 1.1250 ;
        RECT 4.8825 0.7725 4.9875 1.1250 ;
        RECT 4.7775 0.9750 4.8825 1.1250 ;
        RECT 4.6725 0.7725 4.7775 1.1250 ;
        RECT 4.5675 0.9750 4.6725 1.1250 ;
        RECT 4.4625 0.7725 4.5675 1.1250 ;
        RECT 4.3575 0.9750 4.4625 1.1250 ;
        RECT 4.2525 0.7725 4.3575 1.1250 ;
        RECT 4.1475 0.9750 4.2525 1.1250 ;
        RECT 4.0425 0.7725 4.1475 1.1250 ;
        RECT 3.9375 0.9750 4.0425 1.1250 ;
        RECT 3.8325 0.7725 3.9375 1.1250 ;
        RECT 3.7275 0.9750 3.8325 1.1250 ;
        RECT 3.6225 0.7725 3.7275 1.1250 ;
        RECT 3.5175 0.9750 3.6225 1.1250 ;
        RECT 3.4125 0.7725 3.5175 1.1250 ;
        RECT 3.3075 0.9750 3.4125 1.1250 ;
        RECT 3.2025 0.7725 3.3075 1.1250 ;
        RECT 3.0975 0.9750 3.2025 1.1250 ;
        RECT 2.9925 0.7725 3.0975 1.1250 ;
        RECT 2.8875 0.9750 2.9925 1.1250 ;
        RECT 2.7825 0.7725 2.8875 1.1250 ;
        RECT 2.6775 0.9750 2.7825 1.1250 ;
        RECT 2.5725 0.7725 2.6775 1.1250 ;
        RECT 2.4675 0.9750 2.5725 1.1250 ;
        RECT 2.3625 0.7725 2.4675 1.1250 ;
        RECT 2.2575 0.9750 2.3625 1.1250 ;
        RECT 2.1525 0.7725 2.2575 1.1250 ;
        RECT 2.0475 0.9750 2.1525 1.1250 ;
        RECT 1.9425 0.7725 2.0475 1.1250 ;
        RECT 1.8375 0.9750 1.9425 1.1250 ;
        RECT 1.7325 0.7725 1.8375 1.1250 ;
        RECT 1.6275 0.9750 1.7325 1.1250 ;
        RECT 1.5225 0.7725 1.6275 1.1250 ;
        RECT 1.4175 0.9750 1.5225 1.1250 ;
        RECT 1.3125 0.7725 1.4175 1.1250 ;
        RECT 1.2075 0.9750 1.3125 1.1250 ;
        RECT 1.1025 0.7725 1.2075 1.1250 ;
        RECT 0.9975 0.9750 1.1025 1.1250 ;
        RECT 0.8925 0.7725 0.9975 1.1250 ;
        RECT 0.7875 0.9750 0.8925 1.1250 ;
        RECT 0.6825 0.7725 0.7875 1.1250 ;
        RECT 0.5775 0.9750 0.6825 1.1250 ;
        RECT 0.4725 0.7725 0.5775 1.1250 ;
        RECT 0.3675 0.9750 0.4725 1.1250 ;
        RECT 0.2625 0.7725 0.3675 1.1250 ;
        RECT 0.1575 0.9750 0.2625 1.1250 ;
        RECT 0.0525 0.7725 0.1575 1.1250 ;
        RECT 0.0000 0.9750 0.0525 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 13.3050 0.8025 13.3650 0.8625 ;
        RECT 13.2000 0.6000 13.2600 0.6600 ;
        RECT 13.0950 0.8025 13.1550 0.8625 ;
        RECT 12.9900 0.5550 13.0500 0.6150 ;
        RECT 12.8850 0.8025 12.9450 0.8625 ;
        RECT 12.7800 0.5550 12.8400 0.6150 ;
        RECT 12.6750 0.8025 12.7350 0.8625 ;
        RECT 12.5700 0.5550 12.6300 0.6150 ;
        RECT 12.4650 0.8025 12.5250 0.8625 ;
        RECT 12.3600 0.5550 12.4200 0.6150 ;
        RECT 12.2550 0.8025 12.3150 0.8625 ;
        RECT 12.1500 0.5550 12.2100 0.6150 ;
        RECT 12.0450 0.8025 12.1050 0.8625 ;
        RECT 11.9400 0.5550 12.0000 0.6150 ;
        RECT 11.8350 0.8025 11.8950 0.8625 ;
        RECT 11.7300 0.5550 11.7900 0.6150 ;
        RECT 11.6250 0.8025 11.6850 0.8625 ;
        RECT 11.5200 0.5550 11.5800 0.6150 ;
        RECT 11.4150 0.8025 11.4750 0.8625 ;
        RECT 11.3100 0.5550 11.3700 0.6150 ;
        RECT 11.2050 0.8025 11.2650 0.8625 ;
        RECT 11.1000 0.5550 11.1600 0.6150 ;
        RECT 10.9950 0.8025 11.0550 0.8625 ;
        RECT 10.8900 0.5550 10.9500 0.6150 ;
        RECT 10.7850 0.8025 10.8450 0.8625 ;
        RECT 10.6800 0.5550 10.7400 0.6150 ;
        RECT 10.5750 0.8025 10.6350 0.8625 ;
        RECT 10.4700 0.5550 10.5300 0.6150 ;
        RECT 10.3650 0.8025 10.4250 0.8625 ;
        RECT 10.2600 0.5550 10.3200 0.6150 ;
        RECT 10.1550 0.8025 10.2150 0.8625 ;
        RECT 10.0500 0.5550 10.1100 0.6150 ;
        RECT 9.9450 0.8025 10.0050 0.8625 ;
        RECT 9.8400 0.5550 9.9000 0.6150 ;
        RECT 9.7350 0.8025 9.7950 0.8625 ;
        RECT 9.6300 0.5550 9.6900 0.6150 ;
        RECT 9.5250 0.8025 9.5850 0.8625 ;
        RECT 9.4200 0.5550 9.4800 0.6150 ;
        RECT 9.3150 0.8025 9.3750 0.8625 ;
        RECT 9.2100 0.5550 9.2700 0.6150 ;
        RECT 9.1050 0.8025 9.1650 0.8625 ;
        RECT 9.0000 0.5550 9.0600 0.6150 ;
        RECT 8.8950 0.8025 8.9550 0.8625 ;
        RECT 8.7900 0.5550 8.8500 0.6150 ;
        RECT 8.6850 0.8025 8.7450 0.8625 ;
        RECT 8.5800 0.5550 8.6400 0.6150 ;
        RECT 8.4750 0.8025 8.5350 0.8625 ;
        RECT 8.3700 0.5550 8.4300 0.6150 ;
        RECT 8.2650 0.8025 8.3250 0.8625 ;
        RECT 8.1600 0.5550 8.2200 0.6150 ;
        RECT 8.0550 0.8025 8.1150 0.8625 ;
        RECT 7.9500 0.5550 8.0100 0.6150 ;
        RECT 7.8450 0.8025 7.9050 0.8625 ;
        RECT 7.7400 0.5550 7.8000 0.6150 ;
        RECT 7.6350 0.8025 7.6950 0.8625 ;
        RECT 7.5300 0.5550 7.5900 0.6150 ;
        RECT 7.4250 0.8025 7.4850 0.8625 ;
        RECT 7.3200 0.5550 7.3800 0.6150 ;
        RECT 7.2150 0.8025 7.2750 0.8625 ;
        RECT 7.1100 0.5550 7.1700 0.6150 ;
        RECT 7.0050 0.8175 7.0650 0.8775 ;
        RECT 6.7950 0.1875 6.8550 0.2475 ;
        RECT 6.7950 0.8175 6.8550 0.8775 ;
        RECT 6.6900 0.3750 6.7500 0.4350 ;
        RECT 6.6900 0.6150 6.7500 0.6750 ;
        RECT 6.5850 0.1725 6.6450 0.2325 ;
        RECT 6.5850 0.8175 6.6450 0.8775 ;
        RECT 6.4800 0.3750 6.5400 0.4350 ;
        RECT 6.3750 0.1950 6.4350 0.2550 ;
        RECT 6.3750 0.8025 6.4350 0.8625 ;
        RECT 6.2700 0.5550 6.3300 0.6150 ;
        RECT 6.1650 0.8025 6.2250 0.8625 ;
        RECT 6.0600 0.5550 6.1200 0.6150 ;
        RECT 5.9550 0.8025 6.0150 0.8625 ;
        RECT 5.8500 0.5550 5.9100 0.6150 ;
        RECT 5.7450 0.8025 5.8050 0.8625 ;
        RECT 5.6400 0.5550 5.7000 0.6150 ;
        RECT 5.5350 0.8025 5.5950 0.8625 ;
        RECT 5.4300 0.5550 5.4900 0.6150 ;
        RECT 5.3250 0.8025 5.3850 0.8625 ;
        RECT 5.2200 0.5550 5.2800 0.6150 ;
        RECT 5.1150 0.8025 5.1750 0.8625 ;
        RECT 5.0100 0.5550 5.0700 0.6150 ;
        RECT 4.9050 0.8025 4.9650 0.8625 ;
        RECT 4.8000 0.5550 4.8600 0.6150 ;
        RECT 4.6950 0.8025 4.7550 0.8625 ;
        RECT 4.5900 0.5550 4.6500 0.6150 ;
        RECT 4.4850 0.8025 4.5450 0.8625 ;
        RECT 4.3800 0.5550 4.4400 0.6150 ;
        RECT 4.2750 0.8025 4.3350 0.8625 ;
        RECT 4.1700 0.5550 4.2300 0.6150 ;
        RECT 4.0650 0.8025 4.1250 0.8625 ;
        RECT 3.9600 0.5550 4.0200 0.6150 ;
        RECT 3.8550 0.8025 3.9150 0.8625 ;
        RECT 3.7500 0.5550 3.8100 0.6150 ;
        RECT 3.6450 0.8025 3.7050 0.8625 ;
        RECT 3.5400 0.5550 3.6000 0.6150 ;
        RECT 3.4350 0.8025 3.4950 0.8625 ;
        RECT 3.3300 0.5550 3.3900 0.6150 ;
        RECT 3.2250 0.8025 3.2850 0.8625 ;
        RECT 3.1200 0.5550 3.1800 0.6150 ;
        RECT 3.0150 0.8025 3.0750 0.8625 ;
        RECT 2.9100 0.5550 2.9700 0.6150 ;
        RECT 2.8050 0.8025 2.8650 0.8625 ;
        RECT 2.7000 0.5550 2.7600 0.6150 ;
        RECT 2.5950 0.8025 2.6550 0.8625 ;
        RECT 2.4900 0.5550 2.5500 0.6150 ;
        RECT 2.3850 0.8025 2.4450 0.8625 ;
        RECT 2.2800 0.5550 2.3400 0.6150 ;
        RECT 2.1750 0.8025 2.2350 0.8625 ;
        RECT 2.0700 0.5550 2.1300 0.6150 ;
        RECT 1.9650 0.8025 2.0250 0.8625 ;
        RECT 1.8600 0.5550 1.9200 0.6150 ;
        RECT 1.7550 0.8025 1.8150 0.8625 ;
        RECT 1.6500 0.5550 1.7100 0.6150 ;
        RECT 1.5450 0.8025 1.6050 0.8625 ;
        RECT 1.4400 0.5550 1.5000 0.6150 ;
        RECT 1.3350 0.8025 1.3950 0.8625 ;
        RECT 1.2300 0.5550 1.2900 0.6150 ;
        RECT 1.1250 0.8025 1.1850 0.8625 ;
        RECT 1.0200 0.5550 1.0800 0.6150 ;
        RECT 0.9150 0.8025 0.9750 0.8625 ;
        RECT 0.8100 0.5550 0.8700 0.6150 ;
        RECT 0.7050 0.8025 0.7650 0.8625 ;
        RECT 0.6000 0.5550 0.6600 0.6150 ;
        RECT 0.4950 0.8025 0.5550 0.8625 ;
        RECT 0.3900 0.5475 0.4500 0.6075 ;
        RECT 0.2850 0.8025 0.3450 0.8625 ;
        RECT 0.1800 0.6000 0.2400 0.6600 ;
        RECT 0.0750 0.8025 0.1350 0.8625 ;
        LAYER M1 ;
        RECT 13.1700 0.5400 13.2900 0.6600 ;
        RECT 7.1475 0.5400 13.1700 0.6150 ;
        RECT 7.0725 0.1650 7.1475 0.6150 ;
        RECT 6.9300 0.7950 7.0875 0.9000 ;
        RECT 6.7725 0.1650 7.0725 0.2700 ;
        RECT 6.8550 0.3675 6.9300 0.9000 ;
        RECT 6.4425 0.3675 6.8550 0.4425 ;
        RECT 6.7725 0.7950 6.8550 0.9000 ;
        RECT 6.6750 0.6150 6.7800 0.7200 ;
        RECT 6.3375 0.6150 6.6750 0.6900 ;
        RECT 6.3375 0.1725 6.4575 0.2850 ;
        RECT 6.2625 0.1725 6.3375 0.6900 ;
        RECT 0.2700 0.5400 6.2625 0.6150 ;
        RECT 0.1500 0.5400 0.2700 0.6600 ;
        LAYER VIA1 ;
        RECT 7.0725 0.4125 7.1475 0.4875 ;
        RECT 6.2625 0.4125 6.3375 0.4875 ;
        LAYER M2 ;
        RECT 6.1875 0.4125 7.2225 0.4875 ;
    END
END DCAP64_0010


MACRO DCAP8_0010
    CLASS CORE ;
    FOREIGN DCAP8_0010 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.6800 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.1575 -0.0750 1.6800 0.0750 ;
        RECT 0.0525 -0.0750 0.1575 0.2625 ;
        RECT 0.0000 -0.0750 0.0525 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.6275 0.9750 1.6800 1.1250 ;
        RECT 1.5225 0.7725 1.6275 1.1250 ;
        RECT 1.4175 0.9750 1.5225 1.1250 ;
        RECT 1.3125 0.7725 1.4175 1.1250 ;
        RECT 1.2075 0.9750 1.3125 1.1250 ;
        RECT 1.1025 0.7725 1.2075 1.1250 ;
        RECT 0.9975 0.9750 1.1025 1.1250 ;
        RECT 0.8925 0.7725 0.9975 1.1250 ;
        RECT 0.7875 0.9750 0.8925 1.1250 ;
        RECT 0.6825 0.7725 0.7875 1.1250 ;
        RECT 0.5625 0.9750 0.6825 1.1250 ;
        RECT 0.4875 0.7725 0.5625 1.1250 ;
        RECT 0.1575 0.9750 0.4875 1.1250 ;
        RECT 0.0525 0.7725 0.1575 1.1250 ;
        RECT 0.0000 0.9750 0.0525 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.5450 0.8025 1.6050 0.8625 ;
        RECT 1.4400 0.6000 1.5000 0.6600 ;
        RECT 1.3350 0.8025 1.3950 0.8625 ;
        RECT 1.2300 0.5475 1.2900 0.6075 ;
        RECT 1.1250 0.8025 1.1850 0.8625 ;
        RECT 1.0200 0.5550 1.0800 0.6150 ;
        RECT 0.9150 0.8025 0.9750 0.8625 ;
        RECT 0.8100 0.5550 0.8700 0.6150 ;
        RECT 0.7050 0.8025 0.7650 0.8625 ;
        RECT 0.6000 0.5550 0.6600 0.6150 ;
        RECT 0.4950 0.8025 0.5550 0.8625 ;
        RECT 0.2850 0.1800 0.3450 0.2400 ;
        RECT 0.2850 0.7950 0.3450 0.8550 ;
        RECT 0.1800 0.3600 0.2400 0.4200 ;
        RECT 0.1800 0.6000 0.2400 0.6600 ;
        RECT 0.0750 0.1725 0.1350 0.2325 ;
        RECT 0.0750 0.8025 0.1350 0.8625 ;
        LAYER M1 ;
        RECT 1.4100 0.5400 1.5300 0.6600 ;
        RECT 0.7125 0.5400 1.4100 0.6150 ;
        RECT 0.6750 0.5400 0.7125 0.6525 ;
        RECT 0.6000 0.1575 0.6750 0.6525 ;
        RECT 0.2625 0.1575 0.6000 0.2625 ;
        RECT 0.5250 0.5400 0.6000 0.6525 ;
        RECT 0.3375 0.3525 0.4125 0.8775 ;
        RECT 0.1275 0.3525 0.3375 0.4275 ;
        RECT 0.2550 0.7725 0.3375 0.8775 ;
        RECT 0.0975 0.5025 0.2625 0.6975 ;
        LAYER VIA1 ;
        RECT 0.5625 0.5625 0.6375 0.6375 ;
        RECT 0.1725 0.5625 0.2475 0.6375 ;
        LAYER M2 ;
        RECT 0.0975 0.5625 0.7125 0.6375 ;
    END
END DCAP8_0010


MACRO DCCKB_0100
    CLASS CORE ;
    FOREIGN DCCKB_0100 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.0400 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 1.7325 0.2625 1.8900 0.3825 ;
        RECT 1.7325 0.6600 1.8900 0.7800 ;
        RECT 1.4175 0.2625 1.7325 0.7800 ;
        RECT 1.2600 0.2625 1.4175 0.3825 ;
        RECT 1.2600 0.6600 1.4175 0.7800 ;
        VIA 1.7325 0.3225 VIA12_slot ;
        VIA 1.7325 0.7200 VIA12_slot ;
        VIA 1.4175 0.3225 VIA12_slot ;
        VIA 1.4175 0.7200 VIA12_slot ;
        END
    END Z
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.6450 0.4125 1.1100 0.4875 ;
        RECT 0.4800 0.4125 0.6450 0.5175 ;
        VIA 0.5625 0.4650 VIA12_square ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 4.3500 -0.0750 5.0400 0.0750 ;
        RECT 4.2525 -0.0750 4.3500 0.2625 ;
        RECT 2.4525 -0.0750 4.2525 0.0750 ;
        RECT 2.3775 -0.0750 2.4525 0.2925 ;
        RECT 2.0550 -0.0750 2.3775 0.0750 ;
        RECT 1.9350 -0.0750 2.0550 0.1875 ;
        RECT 1.6350 -0.0750 1.9350 0.0750 ;
        RECT 1.5150 -0.0750 1.6350 0.1875 ;
        RECT 1.2150 -0.0750 1.5150 0.0750 ;
        RECT 1.0950 -0.0750 1.2150 0.1875 ;
        RECT 0.7950 -0.0750 1.0950 0.0750 ;
        RECT 0.6750 -0.0750 0.7950 0.1875 ;
        RECT 0.3750 -0.0750 0.6750 0.0750 ;
        RECT 0.2550 -0.0750 0.3750 0.1875 ;
        RECT 0.0000 -0.0750 0.2550 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 4.9875 0.9750 5.0400 1.1250 ;
        RECT 4.8825 0.7725 4.9875 1.1250 ;
        RECT 4.7775 0.9750 4.8825 1.1250 ;
        RECT 4.6725 0.7725 4.7775 1.1250 ;
        RECT 4.5675 0.9750 4.6725 1.1250 ;
        RECT 4.4625 0.7725 4.5675 1.1250 ;
        RECT 4.3575 0.9750 4.4625 1.1250 ;
        RECT 4.2525 0.7725 4.3575 1.1250 ;
        RECT 4.1475 0.9750 4.2525 1.1250 ;
        RECT 4.0425 0.7725 4.1475 1.1250 ;
        RECT 3.9375 0.9750 4.0425 1.1250 ;
        RECT 3.8325 0.7725 3.9375 1.1250 ;
        RECT 3.7275 0.9750 3.8325 1.1250 ;
        RECT 3.6225 0.7725 3.7275 1.1250 ;
        RECT 3.5175 0.9750 3.6225 1.1250 ;
        RECT 3.4125 0.7725 3.5175 1.1250 ;
        RECT 3.3075 0.9750 3.4125 1.1250 ;
        RECT 3.2025 0.7725 3.3075 1.1250 ;
        RECT 3.0975 0.9750 3.2025 1.1250 ;
        RECT 2.9925 0.7725 3.0975 1.1250 ;
        RECT 2.8875 0.9750 2.9925 1.1250 ;
        RECT 2.7825 0.7725 2.8875 1.1250 ;
        RECT 2.4525 0.9750 2.7825 1.1250 ;
        RECT 2.3775 0.6375 2.4525 1.1250 ;
        RECT 2.0550 0.9750 2.3775 1.1250 ;
        RECT 1.9350 0.8550 2.0550 1.1250 ;
        RECT 1.6350 0.9750 1.9350 1.1250 ;
        RECT 1.5150 0.8550 1.6350 1.1250 ;
        RECT 1.2150 0.9750 1.5150 1.1250 ;
        RECT 1.0950 0.8550 1.2150 1.1250 ;
        RECT 0.7950 0.9750 1.0950 1.1250 ;
        RECT 0.6750 0.8175 0.7950 1.1250 ;
        RECT 0.3675 0.9750 0.6750 1.1250 ;
        RECT 0.2625 0.8100 0.3675 1.1250 ;
        RECT 0.0000 0.9750 0.2625 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 4.9050 0.8025 4.9650 0.8625 ;
        RECT 4.8000 0.6000 4.8600 0.6600 ;
        RECT 4.6950 0.8025 4.7550 0.8625 ;
        RECT 4.5900 0.6000 4.6500 0.6600 ;
        RECT 4.4850 0.1800 4.5450 0.2400 ;
        RECT 4.4850 0.8025 4.5450 0.8625 ;
        RECT 4.3800 0.3600 4.4400 0.4200 ;
        RECT 4.3800 0.6000 4.4400 0.6600 ;
        RECT 4.2750 0.1725 4.3350 0.2325 ;
        RECT 4.2750 0.8025 4.3350 0.8625 ;
        RECT 4.1700 0.5475 4.2300 0.6075 ;
        RECT 4.0650 0.8025 4.1250 0.8625 ;
        RECT 3.9600 0.5550 4.0200 0.6150 ;
        RECT 3.8550 0.8025 3.9150 0.8625 ;
        RECT 3.7500 0.5550 3.8100 0.6150 ;
        RECT 3.6450 0.8025 3.7050 0.8625 ;
        RECT 3.5400 0.5550 3.6000 0.6150 ;
        RECT 3.4350 0.8025 3.4950 0.8625 ;
        RECT 3.3300 0.5550 3.3900 0.6150 ;
        RECT 3.2250 0.8025 3.2850 0.8625 ;
        RECT 3.1200 0.5550 3.1800 0.6150 ;
        RECT 3.0150 0.8025 3.0750 0.8625 ;
        RECT 2.9100 0.5550 2.9700 0.6150 ;
        RECT 2.8050 0.8025 2.8650 0.8625 ;
        RECT 2.7000 0.5550 2.7600 0.6150 ;
        RECT 2.5950 0.7875 2.6550 0.8475 ;
        RECT 2.3850 0.1875 2.4450 0.2475 ;
        RECT 2.3850 0.6675 2.4450 0.7275 ;
        RECT 2.3850 0.8325 2.4450 0.8925 ;
        RECT 2.2800 0.4650 2.3400 0.5250 ;
        RECT 2.1750 0.2850 2.2350 0.3450 ;
        RECT 2.1750 0.6900 2.2350 0.7500 ;
        RECT 2.0700 0.4650 2.1300 0.5250 ;
        RECT 1.9650 0.1275 2.0250 0.1875 ;
        RECT 1.9650 0.8625 2.0250 0.9225 ;
        RECT 1.8600 0.4650 1.9200 0.5250 ;
        RECT 1.7550 0.2850 1.8150 0.3450 ;
        RECT 1.7550 0.6900 1.8150 0.7500 ;
        RECT 1.6500 0.4650 1.7100 0.5250 ;
        RECT 1.5450 0.1275 1.6050 0.1875 ;
        RECT 1.5450 0.8625 1.6050 0.9225 ;
        RECT 1.4400 0.4650 1.5000 0.5250 ;
        RECT 1.3350 0.2850 1.3950 0.3450 ;
        RECT 1.3350 0.6900 1.3950 0.7500 ;
        RECT 1.2300 0.4650 1.2900 0.5250 ;
        RECT 1.1250 0.1275 1.1850 0.1875 ;
        RECT 1.1250 0.8625 1.1850 0.9225 ;
        RECT 1.0200 0.4650 1.0800 0.5250 ;
        RECT 0.9150 0.2850 0.9750 0.3450 ;
        RECT 0.9150 0.6900 0.9750 0.7500 ;
        RECT 0.8100 0.4650 0.8700 0.5250 ;
        RECT 0.7050 0.1275 0.7650 0.1875 ;
        RECT 0.7050 0.8250 0.7650 0.8850 ;
        RECT 0.6000 0.4650 0.6600 0.5250 ;
        RECT 0.4950 0.2700 0.5550 0.3300 ;
        RECT 0.4950 0.6675 0.5550 0.7275 ;
        RECT 0.3900 0.4650 0.4500 0.5250 ;
        RECT 0.2850 0.1275 0.3450 0.1875 ;
        RECT 0.2850 0.8325 0.3450 0.8925 ;
        RECT 0.1800 0.4650 0.2400 0.5250 ;
        RECT 0.0750 0.2250 0.1350 0.2850 ;
        RECT 0.0750 0.7575 0.1350 0.8175 ;
        LAYER M1 ;
        RECT 4.6500 0.5850 4.9050 0.6675 ;
        RECT 4.5750 0.1725 4.6500 0.6675 ;
        RECT 4.4550 0.1725 4.5750 0.2475 ;
        RECT 4.2600 0.5775 4.5750 0.6675 ;
        RECT 2.6250 0.3525 4.4700 0.4275 ;
        RECT 4.1475 0.5400 4.2600 0.6675 ;
        RECT 2.8050 0.5400 4.1475 0.6150 ;
        RECT 2.7000 0.5250 2.8050 0.6450 ;
        RECT 2.6250 0.7575 2.6625 0.8850 ;
        RECT 2.5500 0.3525 2.6250 0.8850 ;
        RECT 0.8175 0.4575 2.3700 0.5325 ;
        RECT 0.8925 0.2625 2.2575 0.3825 ;
        RECT 0.8925 0.6600 2.2575 0.7800 ;
        RECT 0.7425 0.2625 0.8175 0.7350 ;
        RECT 0.1575 0.2625 0.7425 0.3375 ;
        RECT 0.1425 0.6600 0.7425 0.7350 ;
        RECT 0.1125 0.4275 0.6600 0.5625 ;
        RECT 0.0525 0.1950 0.1575 0.3375 ;
        RECT 0.0675 0.6600 0.1425 0.8700 ;
        LAYER M2 ;
        RECT 1.7625 0.2625 1.8900 0.3825 ;
        RECT 1.7625 0.6600 1.8900 0.7800 ;
        RECT 1.2600 0.2625 1.3875 0.3825 ;
        RECT 1.2600 0.6600 1.3875 0.7800 ;
    END
END DCCKB_0100


MACRO DCCKB_0101
    CLASS CORE ;
    FOREIGN DCCKB_0101 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.1400 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 2.3625 0.2625 2.5200 0.3825 ;
        RECT 2.3625 0.6600 2.5200 0.7800 ;
        RECT 2.0475 0.2625 2.3625 0.7800 ;
        RECT 1.8900 0.2625 2.0475 0.3825 ;
        RECT 1.8900 0.6600 2.0475 0.7800 ;
        VIA 2.3625 0.3225 VIA12_slot ;
        VIA 2.3625 0.7200 VIA12_slot ;
        VIA 2.0475 0.3225 VIA12_slot ;
        VIA 2.0475 0.7200 VIA12_slot ;
        END
    END Z
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1425 0.4275 0.8700 0.5625 ;
        RECT 0.0675 0.3675 0.1425 0.6825 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 5.1900 -0.0750 7.1400 0.0750 ;
        RECT 5.0850 -0.0750 5.1900 0.2475 ;
        RECT 3.5250 -0.0750 5.0850 0.0750 ;
        RECT 3.4050 -0.0750 3.5250 0.2925 ;
        RECT 3.1050 -0.0750 3.4050 0.0750 ;
        RECT 2.9850 -0.0750 3.1050 0.1875 ;
        RECT 2.6850 -0.0750 2.9850 0.0750 ;
        RECT 2.5650 -0.0750 2.6850 0.1875 ;
        RECT 2.2650 -0.0750 2.5650 0.0750 ;
        RECT 2.1450 -0.0750 2.2650 0.1875 ;
        RECT 1.8450 -0.0750 2.1450 0.0750 ;
        RECT 1.7250 -0.0750 1.8450 0.1875 ;
        RECT 1.4250 -0.0750 1.7250 0.0750 ;
        RECT 1.3050 -0.0750 1.4250 0.1875 ;
        RECT 1.0050 -0.0750 1.3050 0.0750 ;
        RECT 0.8850 -0.0750 1.0050 0.1875 ;
        RECT 0.5850 -0.0750 0.8850 0.0750 ;
        RECT 0.4650 -0.0750 0.5850 0.1875 ;
        RECT 0.1575 -0.0750 0.4650 0.0750 ;
        RECT 0.0525 -0.0750 0.1575 0.2475 ;
        RECT 0.0000 -0.0750 0.0525 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 7.0875 0.9750 7.1400 1.1250 ;
        RECT 6.9825 0.7725 7.0875 1.1250 ;
        RECT 6.8775 0.9750 6.9825 1.1250 ;
        RECT 6.7725 0.7725 6.8775 1.1250 ;
        RECT 6.6675 0.9750 6.7725 1.1250 ;
        RECT 6.5625 0.7725 6.6675 1.1250 ;
        RECT 6.4575 0.9750 6.5625 1.1250 ;
        RECT 6.3525 0.7725 6.4575 1.1250 ;
        RECT 6.2475 0.9750 6.3525 1.1250 ;
        RECT 6.1425 0.7725 6.2475 1.1250 ;
        RECT 6.0375 0.9750 6.1425 1.1250 ;
        RECT 5.9325 0.7725 6.0375 1.1250 ;
        RECT 5.8275 0.9750 5.9325 1.1250 ;
        RECT 5.7225 0.7725 5.8275 1.1250 ;
        RECT 5.6175 0.9750 5.7225 1.1250 ;
        RECT 5.5125 0.7725 5.6175 1.1250 ;
        RECT 5.4075 0.9750 5.5125 1.1250 ;
        RECT 5.3025 0.7725 5.4075 1.1250 ;
        RECT 5.1975 0.9750 5.3025 1.1250 ;
        RECT 5.0925 0.7725 5.1975 1.1250 ;
        RECT 4.9875 0.9750 5.0925 1.1250 ;
        RECT 4.8825 0.7725 4.9875 1.1250 ;
        RECT 4.7775 0.9750 4.8825 1.1250 ;
        RECT 4.6725 0.7725 4.7775 1.1250 ;
        RECT 4.5675 0.9750 4.6725 1.1250 ;
        RECT 4.4625 0.7725 4.5675 1.1250 ;
        RECT 4.3575 0.9750 4.4625 1.1250 ;
        RECT 4.2525 0.7725 4.3575 1.1250 ;
        RECT 4.1475 0.9750 4.2525 1.1250 ;
        RECT 4.0425 0.7725 4.1475 1.1250 ;
        RECT 3.9375 0.9750 4.0425 1.1250 ;
        RECT 3.8325 0.7725 3.9375 1.1250 ;
        RECT 3.5250 0.9750 3.8325 1.1250 ;
        RECT 3.4050 0.6375 3.5250 1.1250 ;
        RECT 3.1050 0.9750 3.4050 1.1250 ;
        RECT 2.9850 0.8550 3.1050 1.1250 ;
        RECT 2.6850 0.9750 2.9850 1.1250 ;
        RECT 2.5650 0.8550 2.6850 1.1250 ;
        RECT 2.2650 0.9750 2.5650 1.1250 ;
        RECT 2.1450 0.8550 2.2650 1.1250 ;
        RECT 1.8450 0.9750 2.1450 1.1250 ;
        RECT 1.7250 0.8550 1.8450 1.1250 ;
        RECT 1.4250 0.9750 1.7250 1.1250 ;
        RECT 1.3050 0.8550 1.4250 1.1250 ;
        RECT 1.0050 0.9750 1.3050 1.1250 ;
        RECT 0.8850 0.8175 1.0050 1.1250 ;
        RECT 0.5775 0.9750 0.8850 1.1250 ;
        RECT 0.4725 0.8100 0.5775 1.1250 ;
        RECT 0.1575 0.9750 0.4725 1.1250 ;
        RECT 0.0525 0.8025 0.1575 1.1250 ;
        RECT 0.0000 0.9750 0.0525 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 7.0050 0.8025 7.0650 0.8625 ;
        RECT 6.9000 0.5550 6.9600 0.6150 ;
        RECT 6.7950 0.8025 6.8550 0.8625 ;
        RECT 6.6900 0.5550 6.7500 0.6150 ;
        RECT 6.5850 0.8025 6.6450 0.8625 ;
        RECT 6.4800 0.5550 6.5400 0.6150 ;
        RECT 6.3750 0.8025 6.4350 0.8625 ;
        RECT 6.2700 0.5550 6.3300 0.6150 ;
        RECT 6.1650 0.8025 6.2250 0.8625 ;
        RECT 6.0600 0.5550 6.1200 0.6150 ;
        RECT 5.9550 0.8025 6.0150 0.8625 ;
        RECT 5.8500 0.5550 5.9100 0.6150 ;
        RECT 5.7450 0.8025 5.8050 0.8625 ;
        RECT 5.6400 0.5550 5.7000 0.6150 ;
        RECT 5.5350 0.8025 5.5950 0.8625 ;
        RECT 5.4300 0.5475 5.4900 0.6075 ;
        RECT 5.3250 0.1575 5.3850 0.2175 ;
        RECT 5.3250 0.8025 5.3850 0.8625 ;
        RECT 5.2200 0.3300 5.2800 0.3900 ;
        RECT 5.2200 0.5700 5.2800 0.6300 ;
        RECT 5.1150 0.1575 5.1750 0.2175 ;
        RECT 5.1150 0.8025 5.1750 0.8625 ;
        RECT 5.0100 0.5475 5.0700 0.6075 ;
        RECT 4.9050 0.8025 4.9650 0.8625 ;
        RECT 4.8000 0.5550 4.8600 0.6150 ;
        RECT 4.6950 0.8025 4.7550 0.8625 ;
        RECT 4.5900 0.5550 4.6500 0.6150 ;
        RECT 4.4850 0.8025 4.5450 0.8625 ;
        RECT 4.3800 0.5550 4.4400 0.6150 ;
        RECT 4.2750 0.8025 4.3350 0.8625 ;
        RECT 4.1700 0.5550 4.2300 0.6150 ;
        RECT 4.0650 0.8025 4.1250 0.8625 ;
        RECT 3.9600 0.5550 4.0200 0.6150 ;
        RECT 3.8550 0.8025 3.9150 0.8625 ;
        RECT 3.7500 0.5550 3.8100 0.6150 ;
        RECT 3.6450 0.7875 3.7050 0.8475 ;
        RECT 3.4350 0.1875 3.4950 0.2475 ;
        RECT 3.4350 0.6675 3.4950 0.7275 ;
        RECT 3.4350 0.8325 3.4950 0.8925 ;
        RECT 3.3300 0.4650 3.3900 0.5250 ;
        RECT 3.2250 0.2925 3.2850 0.3525 ;
        RECT 3.2250 0.6900 3.2850 0.7500 ;
        RECT 3.1200 0.4650 3.1800 0.5250 ;
        RECT 3.0150 0.1275 3.0750 0.1875 ;
        RECT 3.0150 0.8625 3.0750 0.9225 ;
        RECT 2.9100 0.4650 2.9700 0.5250 ;
        RECT 2.8050 0.2925 2.8650 0.3525 ;
        RECT 2.8050 0.6900 2.8650 0.7500 ;
        RECT 2.7000 0.4650 2.7600 0.5250 ;
        RECT 2.5950 0.1275 2.6550 0.1875 ;
        RECT 2.5950 0.8625 2.6550 0.9225 ;
        RECT 2.4900 0.4650 2.5500 0.5250 ;
        RECT 2.3850 0.2925 2.4450 0.3525 ;
        RECT 2.3850 0.6900 2.4450 0.7500 ;
        RECT 2.2800 0.4650 2.3400 0.5250 ;
        RECT 2.1750 0.1275 2.2350 0.1875 ;
        RECT 2.1750 0.8625 2.2350 0.9225 ;
        RECT 2.0700 0.4650 2.1300 0.5250 ;
        RECT 1.9650 0.2925 2.0250 0.3525 ;
        RECT 1.9650 0.6900 2.0250 0.7500 ;
        RECT 1.8600 0.4650 1.9200 0.5250 ;
        RECT 1.7550 0.1275 1.8150 0.1875 ;
        RECT 1.7550 0.8625 1.8150 0.9225 ;
        RECT 1.6500 0.4650 1.7100 0.5250 ;
        RECT 1.5450 0.2925 1.6050 0.3525 ;
        RECT 1.5450 0.6900 1.6050 0.7500 ;
        RECT 1.4400 0.4650 1.5000 0.5250 ;
        RECT 1.3350 0.1275 1.3950 0.1875 ;
        RECT 1.3350 0.8625 1.3950 0.9225 ;
        RECT 1.2300 0.4650 1.2900 0.5250 ;
        RECT 1.1250 0.2925 1.1850 0.3525 ;
        RECT 1.1250 0.6900 1.1850 0.7500 ;
        RECT 1.0200 0.4650 1.0800 0.5250 ;
        RECT 0.9150 0.1275 0.9750 0.1875 ;
        RECT 0.9150 0.8250 0.9750 0.8850 ;
        RECT 0.8100 0.4650 0.8700 0.5250 ;
        RECT 0.7050 0.2700 0.7650 0.3300 ;
        RECT 0.7050 0.6675 0.7650 0.7275 ;
        RECT 0.6000 0.4650 0.6600 0.5250 ;
        RECT 0.4950 0.1275 0.5550 0.1875 ;
        RECT 0.4950 0.8325 0.5550 0.8925 ;
        RECT 0.3900 0.4650 0.4500 0.5250 ;
        RECT 0.2850 0.2250 0.3450 0.2850 ;
        RECT 0.2850 0.7050 0.3450 0.7650 ;
        RECT 0.1800 0.4650 0.2400 0.5250 ;
        RECT 0.0750 0.1575 0.1350 0.2175 ;
        RECT 0.0750 0.8325 0.1350 0.8925 ;
        LAYER M1 ;
        RECT 5.4600 0.5475 7.0050 0.6300 ;
        RECT 5.3850 0.1500 5.4600 0.6300 ;
        RECT 5.2950 0.1500 5.3850 0.2250 ;
        RECT 3.8550 0.5400 5.3850 0.6300 ;
        RECT 5.1900 0.3225 5.3100 0.4275 ;
        RECT 3.6750 0.3225 5.1900 0.3975 ;
        RECT 3.7500 0.5175 3.8550 0.6450 ;
        RECT 3.6750 0.7575 3.7125 0.8850 ;
        RECT 3.6000 0.3225 3.6750 0.8850 ;
        RECT 1.0275 0.4575 3.4200 0.5325 ;
        RECT 1.1025 0.2625 3.3075 0.3825 ;
        RECT 1.1025 0.6600 3.3075 0.7800 ;
        RECT 0.9525 0.2625 1.0275 0.7350 ;
        RECT 0.3525 0.2625 0.9525 0.3375 ;
        RECT 0.3525 0.6600 0.9525 0.7350 ;
        RECT 0.2775 0.1950 0.3525 0.3375 ;
        RECT 0.2775 0.6600 0.3525 0.8100 ;
        LAYER M2 ;
        RECT 2.3925 0.2625 2.5200 0.3825 ;
        RECT 2.3925 0.6600 2.5200 0.7800 ;
        RECT 1.8900 0.2625 2.0175 0.3825 ;
        RECT 1.8900 0.6600 2.0175 0.7800 ;
    END
END DCCKB_0101


MACRO DCCKB_0111
    CLASS CORE ;
    FOREIGN DCCKB_0111 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.9400 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 0.7875 0.2625 1.1025 0.7500 ;
        VIA 0.9450 0.3450 VIA12_slot ;
        VIA 0.9450 0.6675 VIA12_slot ;
        END
    END Z
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1575 0.4275 0.4500 0.5625 ;
        RECT 0.0525 0.3675 0.1575 0.6825 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 2.2500 -0.0750 2.9400 0.0750 ;
        RECT 2.1525 -0.0750 2.2500 0.2625 ;
        RECT 1.4025 -0.0750 2.1525 0.0750 ;
        RECT 1.3275 -0.0750 1.4025 0.3150 ;
        RECT 1.0050 -0.0750 1.3275 0.0750 ;
        RECT 0.8850 -0.0750 1.0050 0.1950 ;
        RECT 0.5850 -0.0750 0.8850 0.0750 ;
        RECT 0.4650 -0.0750 0.5850 0.1875 ;
        RECT 0.1425 -0.0750 0.4650 0.0750 ;
        RECT 0.0675 -0.0750 0.1425 0.2625 ;
        RECT 0.0000 -0.0750 0.0675 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 2.8875 0.9750 2.9400 1.1250 ;
        RECT 2.7825 0.7725 2.8875 1.1250 ;
        RECT 2.6775 0.9750 2.7825 1.1250 ;
        RECT 2.5725 0.7725 2.6775 1.1250 ;
        RECT 2.4675 0.9750 2.5725 1.1250 ;
        RECT 2.3625 0.7725 2.4675 1.1250 ;
        RECT 2.2575 0.9750 2.3625 1.1250 ;
        RECT 2.1525 0.7725 2.2575 1.1250 ;
        RECT 2.0475 0.9750 2.1525 1.1250 ;
        RECT 1.9425 0.7725 2.0475 1.1250 ;
        RECT 1.8375 0.9750 1.9425 1.1250 ;
        RECT 1.7325 0.7725 1.8375 1.1250 ;
        RECT 1.4175 0.9750 1.7325 1.1250 ;
        RECT 1.3125 0.6375 1.4175 1.1250 ;
        RECT 0.9825 0.9750 1.3125 1.1250 ;
        RECT 0.9075 0.8175 0.9825 1.1250 ;
        RECT 0.5850 0.9750 0.9075 1.1250 ;
        RECT 0.4650 0.8175 0.5850 1.1250 ;
        RECT 0.1425 0.9750 0.4650 1.1250 ;
        RECT 0.0675 0.7950 0.1425 1.1250 ;
        RECT 0.0000 0.9750 0.0675 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 2.8050 0.8025 2.8650 0.8625 ;
        RECT 2.7000 0.6000 2.7600 0.6600 ;
        RECT 2.5950 0.8025 2.6550 0.8625 ;
        RECT 2.4900 0.6000 2.5500 0.6600 ;
        RECT 2.3850 0.1800 2.4450 0.2400 ;
        RECT 2.3850 0.8025 2.4450 0.8625 ;
        RECT 2.2800 0.3600 2.3400 0.4200 ;
        RECT 2.2800 0.6000 2.3400 0.6600 ;
        RECT 2.1750 0.1725 2.2350 0.2325 ;
        RECT 2.1750 0.8025 2.2350 0.8625 ;
        RECT 2.0700 0.5475 2.1300 0.6075 ;
        RECT 1.9650 0.8025 2.0250 0.8625 ;
        RECT 1.8600 0.5550 1.9200 0.6150 ;
        RECT 1.7550 0.8025 1.8150 0.8625 ;
        RECT 1.6500 0.5550 1.7100 0.6150 ;
        RECT 1.5450 0.7875 1.6050 0.8475 ;
        RECT 1.3350 0.2250 1.3950 0.2850 ;
        RECT 1.3350 0.6675 1.3950 0.7275 ;
        RECT 1.3350 0.8325 1.3950 0.8925 ;
        RECT 1.2300 0.4800 1.2900 0.5400 ;
        RECT 1.1250 0.2250 1.1850 0.2850 ;
        RECT 1.1250 0.7575 1.1850 0.8175 ;
        RECT 1.0200 0.4800 1.0800 0.5400 ;
        RECT 0.9150 0.1275 0.9750 0.1875 ;
        RECT 0.9150 0.8475 0.9750 0.9075 ;
        RECT 0.8100 0.4800 0.8700 0.5400 ;
        RECT 0.7050 0.2250 0.7650 0.2850 ;
        RECT 0.7050 0.7575 0.7650 0.8175 ;
        RECT 0.6000 0.4800 0.6600 0.5400 ;
        RECT 0.4950 0.1275 0.5550 0.1875 ;
        RECT 0.4950 0.8250 0.5550 0.8850 ;
        RECT 0.3900 0.4650 0.4500 0.5250 ;
        RECT 0.2850 0.2250 0.3450 0.2850 ;
        RECT 0.2850 0.7575 0.3450 0.8175 ;
        RECT 0.1800 0.4650 0.2400 0.5250 ;
        RECT 0.0750 0.1725 0.1350 0.2325 ;
        RECT 0.0750 0.8250 0.1350 0.8850 ;
        LAYER M1 ;
        RECT 2.5500 0.5850 2.8050 0.6675 ;
        RECT 2.4750 0.1725 2.5500 0.6675 ;
        RECT 2.3550 0.1725 2.4750 0.2475 ;
        RECT 2.1600 0.5775 2.4750 0.6675 ;
        RECT 1.5750 0.3525 2.3700 0.4275 ;
        RECT 2.0475 0.5400 2.1600 0.6675 ;
        RECT 1.7550 0.5400 2.0475 0.6150 ;
        RECT 1.6500 0.5250 1.7550 0.6450 ;
        RECT 1.5750 0.7575 1.6125 0.8850 ;
        RECT 1.5000 0.3525 1.5750 0.8850 ;
        RECT 0.6075 0.4725 1.3200 0.5475 ;
        RECT 1.1025 0.1950 1.2075 0.3900 ;
        RECT 1.1175 0.6225 1.1925 0.8700 ;
        RECT 0.7725 0.6225 1.1175 0.7125 ;
        RECT 0.7875 0.3000 1.1025 0.3900 ;
        RECT 0.6825 0.1950 0.7875 0.3900 ;
        RECT 0.6975 0.6225 0.7725 0.8700 ;
        RECT 0.5325 0.2625 0.6075 0.7125 ;
        RECT 0.3675 0.2625 0.5325 0.3375 ;
        RECT 0.3525 0.6375 0.5325 0.7125 ;
        RECT 0.2625 0.1950 0.3675 0.3375 ;
        RECT 0.2775 0.6375 0.3525 0.8700 ;
    END
END DCCKB_0111


MACRO DCCKB_1100
    CLASS CORE ;
    FOREIGN DCCKB_1100 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.2400 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 2.9925 0.2625 3.1500 0.3825 ;
        RECT 2.9925 0.6600 3.1500 0.7800 ;
        RECT 2.6775 0.2625 2.9925 0.7800 ;
        RECT 2.5200 0.2625 2.6775 0.3825 ;
        RECT 2.5200 0.6600 2.6775 0.7800 ;
        VIA 2.9925 0.3225 VIA12_slot ;
        VIA 2.9925 0.7200 VIA12_slot ;
        VIA 2.6775 0.3225 VIA12_slot ;
        VIA 2.6775 0.7200 VIA12_slot ;
        END
    END Z
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.0425 0.4125 1.5300 0.4875 ;
        RECT 0.8775 0.4125 1.0425 0.5175 ;
        VIA 0.9600 0.4650 VIA12_square ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 8.5500 -0.0750 9.2400 0.0750 ;
        RECT 8.4525 -0.0750 8.5500 0.2625 ;
        RECT 4.5525 -0.0750 8.4525 0.0750 ;
        RECT 4.4775 -0.0750 4.5525 0.2925 ;
        RECT 4.1550 -0.0750 4.4775 0.0750 ;
        RECT 4.0350 -0.0750 4.1550 0.1875 ;
        RECT 3.7350 -0.0750 4.0350 0.0750 ;
        RECT 3.6150 -0.0750 3.7350 0.1875 ;
        RECT 3.3150 -0.0750 3.6150 0.0750 ;
        RECT 3.1950 -0.0750 3.3150 0.1875 ;
        RECT 2.8950 -0.0750 3.1950 0.0750 ;
        RECT 2.7750 -0.0750 2.8950 0.1875 ;
        RECT 2.4750 -0.0750 2.7750 0.0750 ;
        RECT 2.3550 -0.0750 2.4750 0.1875 ;
        RECT 2.0550 -0.0750 2.3550 0.0750 ;
        RECT 1.9350 -0.0750 2.0550 0.1875 ;
        RECT 1.6350 -0.0750 1.9350 0.0750 ;
        RECT 1.5150 -0.0750 1.6350 0.1875 ;
        RECT 1.2150 -0.0750 1.5150 0.0750 ;
        RECT 1.0950 -0.0750 1.2150 0.1875 ;
        RECT 0.7950 -0.0750 1.0950 0.0750 ;
        RECT 0.6750 -0.0750 0.7950 0.1875 ;
        RECT 0.3750 -0.0750 0.6750 0.0750 ;
        RECT 0.2550 -0.0750 0.3750 0.1875 ;
        RECT 0.0000 -0.0750 0.2550 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 9.1875 0.9750 9.2400 1.1250 ;
        RECT 9.0825 0.7725 9.1875 1.1250 ;
        RECT 8.9775 0.9750 9.0825 1.1250 ;
        RECT 8.8725 0.7725 8.9775 1.1250 ;
        RECT 8.7675 0.9750 8.8725 1.1250 ;
        RECT 8.6625 0.7725 8.7675 1.1250 ;
        RECT 8.5575 0.9750 8.6625 1.1250 ;
        RECT 8.4525 0.7725 8.5575 1.1250 ;
        RECT 8.3475 0.9750 8.4525 1.1250 ;
        RECT 8.2425 0.7725 8.3475 1.1250 ;
        RECT 8.1375 0.9750 8.2425 1.1250 ;
        RECT 8.0325 0.7725 8.1375 1.1250 ;
        RECT 7.9275 0.9750 8.0325 1.1250 ;
        RECT 7.8225 0.7725 7.9275 1.1250 ;
        RECT 7.7175 0.9750 7.8225 1.1250 ;
        RECT 7.6125 0.7725 7.7175 1.1250 ;
        RECT 7.5075 0.9750 7.6125 1.1250 ;
        RECT 7.4025 0.7725 7.5075 1.1250 ;
        RECT 7.2975 0.9750 7.4025 1.1250 ;
        RECT 7.1925 0.7725 7.2975 1.1250 ;
        RECT 7.0875 0.9750 7.1925 1.1250 ;
        RECT 6.9825 0.7725 7.0875 1.1250 ;
        RECT 6.8775 0.9750 6.9825 1.1250 ;
        RECT 6.7725 0.7725 6.8775 1.1250 ;
        RECT 6.6675 0.9750 6.7725 1.1250 ;
        RECT 6.5625 0.7725 6.6675 1.1250 ;
        RECT 6.4575 0.9750 6.5625 1.1250 ;
        RECT 6.3525 0.7725 6.4575 1.1250 ;
        RECT 6.2475 0.9750 6.3525 1.1250 ;
        RECT 6.1425 0.7725 6.2475 1.1250 ;
        RECT 6.0375 0.9750 6.1425 1.1250 ;
        RECT 5.9325 0.7725 6.0375 1.1250 ;
        RECT 5.8275 0.9750 5.9325 1.1250 ;
        RECT 5.7225 0.7725 5.8275 1.1250 ;
        RECT 5.6175 0.9750 5.7225 1.1250 ;
        RECT 5.5125 0.7725 5.6175 1.1250 ;
        RECT 5.4075 0.9750 5.5125 1.1250 ;
        RECT 5.3025 0.7725 5.4075 1.1250 ;
        RECT 5.1975 0.9750 5.3025 1.1250 ;
        RECT 5.0925 0.7725 5.1975 1.1250 ;
        RECT 4.9875 0.9750 5.0925 1.1250 ;
        RECT 4.8825 0.7725 4.9875 1.1250 ;
        RECT 4.5525 0.9750 4.8825 1.1250 ;
        RECT 4.4775 0.6375 4.5525 1.1250 ;
        RECT 4.1550 0.9750 4.4775 1.1250 ;
        RECT 4.0350 0.8550 4.1550 1.1250 ;
        RECT 3.7350 0.9750 4.0350 1.1250 ;
        RECT 3.6150 0.8550 3.7350 1.1250 ;
        RECT 3.3150 0.9750 3.6150 1.1250 ;
        RECT 3.1950 0.8550 3.3150 1.1250 ;
        RECT 2.8950 0.9750 3.1950 1.1250 ;
        RECT 2.7750 0.8550 2.8950 1.1250 ;
        RECT 2.4750 0.9750 2.7750 1.1250 ;
        RECT 2.3550 0.8550 2.4750 1.1250 ;
        RECT 2.0550 0.9750 2.3550 1.1250 ;
        RECT 1.9350 0.8550 2.0550 1.1250 ;
        RECT 1.6350 0.9750 1.9350 1.1250 ;
        RECT 1.5150 0.8550 1.6350 1.1250 ;
        RECT 1.2150 0.9750 1.5150 1.1250 ;
        RECT 1.0950 0.8175 1.2150 1.1250 ;
        RECT 0.7950 0.9750 1.0950 1.1250 ;
        RECT 0.6750 0.8175 0.7950 1.1250 ;
        RECT 0.3675 0.9750 0.6750 1.1250 ;
        RECT 0.2625 0.8175 0.3675 1.1250 ;
        RECT 0.0000 0.9750 0.2625 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 9.1050 0.8025 9.1650 0.8625 ;
        RECT 9.0000 0.6000 9.0600 0.6600 ;
        RECT 8.8950 0.8025 8.9550 0.8625 ;
        RECT 8.7900 0.6000 8.8500 0.6600 ;
        RECT 8.6850 0.1800 8.7450 0.2400 ;
        RECT 8.6850 0.8025 8.7450 0.8625 ;
        RECT 8.5800 0.3600 8.6400 0.4200 ;
        RECT 8.5800 0.6000 8.6400 0.6600 ;
        RECT 8.4750 0.1725 8.5350 0.2325 ;
        RECT 8.4750 0.8025 8.5350 0.8625 ;
        RECT 8.3700 0.5475 8.4300 0.6075 ;
        RECT 8.2650 0.8025 8.3250 0.8625 ;
        RECT 8.1600 0.5550 8.2200 0.6150 ;
        RECT 8.0550 0.8025 8.1150 0.8625 ;
        RECT 7.9500 0.5550 8.0100 0.6150 ;
        RECT 7.8450 0.8025 7.9050 0.8625 ;
        RECT 7.7400 0.5550 7.8000 0.6150 ;
        RECT 7.6350 0.8025 7.6950 0.8625 ;
        RECT 7.5300 0.5550 7.5900 0.6150 ;
        RECT 7.4250 0.8025 7.4850 0.8625 ;
        RECT 7.3200 0.5550 7.3800 0.6150 ;
        RECT 7.2150 0.8025 7.2750 0.8625 ;
        RECT 7.1100 0.5550 7.1700 0.6150 ;
        RECT 7.0050 0.8025 7.0650 0.8625 ;
        RECT 6.9000 0.5550 6.9600 0.6150 ;
        RECT 6.7950 0.8025 6.8550 0.8625 ;
        RECT 6.6900 0.5550 6.7500 0.6150 ;
        RECT 6.5850 0.8025 6.6450 0.8625 ;
        RECT 6.4800 0.5550 6.5400 0.6150 ;
        RECT 6.3750 0.8025 6.4350 0.8625 ;
        RECT 6.2700 0.5550 6.3300 0.6150 ;
        RECT 6.1650 0.8025 6.2250 0.8625 ;
        RECT 6.0600 0.5550 6.1200 0.6150 ;
        RECT 5.9550 0.8025 6.0150 0.8625 ;
        RECT 5.8500 0.5550 5.9100 0.6150 ;
        RECT 5.7450 0.8025 5.8050 0.8625 ;
        RECT 5.6400 0.5550 5.7000 0.6150 ;
        RECT 5.5350 0.8025 5.5950 0.8625 ;
        RECT 5.4300 0.5550 5.4900 0.6150 ;
        RECT 5.3250 0.8025 5.3850 0.8625 ;
        RECT 5.2200 0.5550 5.2800 0.6150 ;
        RECT 5.1150 0.8025 5.1750 0.8625 ;
        RECT 5.0100 0.5550 5.0700 0.6150 ;
        RECT 4.9050 0.8025 4.9650 0.8625 ;
        RECT 4.8000 0.5550 4.8600 0.6150 ;
        RECT 4.6950 0.7875 4.7550 0.8475 ;
        RECT 4.4850 0.1875 4.5450 0.2475 ;
        RECT 4.4850 0.6675 4.5450 0.7275 ;
        RECT 4.4850 0.8325 4.5450 0.8925 ;
        RECT 4.3800 0.4650 4.4400 0.5250 ;
        RECT 4.2750 0.2925 4.3350 0.3525 ;
        RECT 4.2750 0.6900 4.3350 0.7500 ;
        RECT 4.1700 0.4650 4.2300 0.5250 ;
        RECT 4.0650 0.1275 4.1250 0.1875 ;
        RECT 4.0650 0.8625 4.1250 0.9225 ;
        RECT 3.9600 0.4650 4.0200 0.5250 ;
        RECT 3.8550 0.2925 3.9150 0.3525 ;
        RECT 3.8550 0.6900 3.9150 0.7500 ;
        RECT 3.7500 0.4650 3.8100 0.5250 ;
        RECT 3.6450 0.1275 3.7050 0.1875 ;
        RECT 3.6450 0.8625 3.7050 0.9225 ;
        RECT 3.5400 0.4650 3.6000 0.5250 ;
        RECT 3.4350 0.2925 3.4950 0.3525 ;
        RECT 3.4350 0.6900 3.4950 0.7500 ;
        RECT 3.3300 0.4650 3.3900 0.5250 ;
        RECT 3.2250 0.1275 3.2850 0.1875 ;
        RECT 3.2250 0.8625 3.2850 0.9225 ;
        RECT 3.1200 0.4650 3.1800 0.5250 ;
        RECT 3.0150 0.2925 3.0750 0.3525 ;
        RECT 3.0150 0.6900 3.0750 0.7500 ;
        RECT 2.9100 0.4650 2.9700 0.5250 ;
        RECT 2.8050 0.1275 2.8650 0.1875 ;
        RECT 2.8050 0.8625 2.8650 0.9225 ;
        RECT 2.7000 0.4650 2.7600 0.5250 ;
        RECT 2.5950 0.2925 2.6550 0.3525 ;
        RECT 2.5950 0.6900 2.6550 0.7500 ;
        RECT 2.4900 0.4650 2.5500 0.5250 ;
        RECT 2.3850 0.1275 2.4450 0.1875 ;
        RECT 2.3850 0.8625 2.4450 0.9225 ;
        RECT 2.2800 0.4650 2.3400 0.5250 ;
        RECT 2.1750 0.2925 2.2350 0.3525 ;
        RECT 2.1750 0.6900 2.2350 0.7500 ;
        RECT 2.0700 0.4650 2.1300 0.5250 ;
        RECT 1.9650 0.1275 2.0250 0.1875 ;
        RECT 1.9650 0.8625 2.0250 0.9225 ;
        RECT 1.8600 0.4650 1.9200 0.5250 ;
        RECT 1.7550 0.2925 1.8150 0.3525 ;
        RECT 1.7550 0.6900 1.8150 0.7500 ;
        RECT 1.6500 0.4650 1.7100 0.5250 ;
        RECT 1.5450 0.1275 1.6050 0.1875 ;
        RECT 1.5450 0.8625 1.6050 0.9225 ;
        RECT 1.4400 0.4650 1.5000 0.5250 ;
        RECT 1.3350 0.2925 1.3950 0.3525 ;
        RECT 1.3350 0.6900 1.3950 0.7500 ;
        RECT 1.2300 0.4650 1.2900 0.5250 ;
        RECT 1.1250 0.1275 1.1850 0.1875 ;
        RECT 1.1250 0.8250 1.1850 0.8850 ;
        RECT 1.0200 0.4650 1.0800 0.5250 ;
        RECT 0.9150 0.2700 0.9750 0.3300 ;
        RECT 0.9150 0.6750 0.9750 0.7350 ;
        RECT 0.8100 0.4650 0.8700 0.5250 ;
        RECT 0.7050 0.1275 0.7650 0.1875 ;
        RECT 0.7050 0.8250 0.7650 0.8850 ;
        RECT 0.6000 0.4650 0.6600 0.5250 ;
        RECT 0.4950 0.2700 0.5550 0.3300 ;
        RECT 0.4950 0.6750 0.5550 0.7350 ;
        RECT 0.3900 0.4650 0.4500 0.5250 ;
        RECT 0.2850 0.1275 0.3450 0.1875 ;
        RECT 0.2850 0.8475 0.3450 0.9075 ;
        RECT 0.1800 0.4650 0.2400 0.5250 ;
        RECT 0.0750 0.2250 0.1350 0.2850 ;
        RECT 0.0750 0.7575 0.1350 0.8175 ;
        LAYER M1 ;
        RECT 8.8500 0.5850 9.1050 0.6675 ;
        RECT 8.7750 0.1725 8.8500 0.6675 ;
        RECT 8.6550 0.1725 8.7750 0.2475 ;
        RECT 8.4600 0.5775 8.7750 0.6675 ;
        RECT 4.7250 0.3525 8.6700 0.4275 ;
        RECT 8.3475 0.5400 8.4600 0.6675 ;
        RECT 4.9050 0.5400 8.3475 0.6150 ;
        RECT 4.8000 0.5250 4.9050 0.6450 ;
        RECT 4.7250 0.7575 4.7625 0.8850 ;
        RECT 4.6500 0.3525 4.7250 0.8850 ;
        RECT 1.2375 0.4575 4.4700 0.5325 ;
        RECT 1.3125 0.2625 4.3575 0.3825 ;
        RECT 1.3125 0.6600 4.3575 0.7800 ;
        RECT 1.1625 0.2625 1.2375 0.7425 ;
        RECT 0.1425 0.2625 1.1625 0.3375 ;
        RECT 0.1425 0.6675 1.1625 0.7425 ;
        RECT 0.1125 0.4275 1.0800 0.5625 ;
        RECT 0.0675 0.1950 0.1425 0.3375 ;
        RECT 0.0675 0.6675 0.1425 0.8700 ;
        LAYER M2 ;
        RECT 3.0225 0.2625 3.1500 0.3825 ;
        RECT 3.0225 0.6600 3.1500 0.7800 ;
        RECT 2.5200 0.2625 2.6475 0.3825 ;
        RECT 2.5200 0.6600 2.6475 0.7800 ;
    END
END DCCKB_1100


MACRO DCCKN_0111
    CLASS CORE ;
    FOREIGN DCCKN_0111 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.1000 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 0.3675 0.2700 0.6825 0.7800 ;
        VIA 0.5250 0.3525 VIA12_slot ;
        VIA 0.5250 0.6975 VIA12_slot ;
        END
    END ZN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1425 0.4725 0.9150 0.5475 ;
        RECT 0.0675 0.3675 0.1425 0.6825 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.2075 -0.0750 2.1000 0.0750 ;
        RECT 1.1025 -0.0750 1.2075 0.2475 ;
        RECT 1.0050 -0.0750 1.1025 0.0750 ;
        RECT 0.8850 -0.0750 1.0050 0.2925 ;
        RECT 0.5850 -0.0750 0.8850 0.0750 ;
        RECT 0.4650 -0.0750 0.5850 0.2025 ;
        RECT 0.1425 -0.0750 0.4650 0.0750 ;
        RECT 0.0675 -0.0750 0.1425 0.2475 ;
        RECT 0.0000 -0.0750 0.0675 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 2.0475 0.9750 2.1000 1.1250 ;
        RECT 1.9425 0.7725 2.0475 1.1250 ;
        RECT 1.8375 0.9750 1.9425 1.1250 ;
        RECT 1.7325 0.7725 1.8375 1.1250 ;
        RECT 1.6275 0.9750 1.7325 1.1250 ;
        RECT 1.5225 0.7725 1.6275 1.1250 ;
        RECT 1.4175 0.9750 1.5225 1.1250 ;
        RECT 1.3125 0.7725 1.4175 1.1250 ;
        RECT 1.0050 0.9750 1.3125 1.1250 ;
        RECT 0.8850 0.6600 1.0050 1.1250 ;
        RECT 0.5850 0.9750 0.8850 1.1250 ;
        RECT 0.4650 0.8475 0.5850 1.1250 ;
        RECT 0.1425 0.9750 0.4650 1.1250 ;
        RECT 0.0675 0.8025 0.1425 1.1250 ;
        RECT 0.0000 0.9750 0.0675 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.9650 0.8025 2.0250 0.8625 ;
        RECT 1.8600 0.6000 1.9200 0.6600 ;
        RECT 1.7550 0.8025 1.8150 0.8625 ;
        RECT 1.6500 0.6000 1.7100 0.6600 ;
        RECT 1.5450 0.8025 1.6050 0.8625 ;
        RECT 1.4400 0.6000 1.5000 0.6600 ;
        RECT 1.3350 0.1725 1.3950 0.2325 ;
        RECT 1.3350 0.8025 1.3950 0.8625 ;
        RECT 1.2300 0.3525 1.2900 0.4125 ;
        RECT 1.2300 0.6000 1.2900 0.6600 ;
        RECT 1.1250 0.1575 1.1850 0.2175 ;
        RECT 1.1250 0.7875 1.1850 0.8475 ;
        RECT 0.9150 0.2175 0.9750 0.2775 ;
        RECT 0.9150 0.6675 0.9750 0.7275 ;
        RECT 0.9150 0.8325 0.9750 0.8925 ;
        RECT 0.8100 0.4800 0.8700 0.5400 ;
        RECT 0.7050 0.2325 0.7650 0.2925 ;
        RECT 0.7050 0.6825 0.7650 0.7425 ;
        RECT 0.6000 0.4800 0.6600 0.5400 ;
        RECT 0.4950 0.1350 0.5550 0.1950 ;
        RECT 0.4950 0.8550 0.5550 0.9150 ;
        RECT 0.3900 0.4800 0.4500 0.5400 ;
        RECT 0.2850 0.2325 0.3450 0.2925 ;
        RECT 0.2850 0.6825 0.3450 0.7425 ;
        RECT 0.1800 0.4800 0.2400 0.5400 ;
        RECT 0.0750 0.1575 0.1350 0.2175 ;
        RECT 0.0750 0.8325 0.1350 0.8925 ;
        LAYER M1 ;
        RECT 1.5450 0.5850 1.9650 0.6750 ;
        RECT 1.4700 0.1500 1.5450 0.6750 ;
        RECT 1.3125 0.1500 1.4700 0.2550 ;
        RECT 1.3350 0.5850 1.4700 0.6750 ;
        RECT 1.2300 0.5700 1.3350 0.6900 ;
        RECT 1.1550 0.3300 1.3125 0.4350 ;
        RECT 1.1550 0.7575 1.1925 0.8850 ;
        RECT 1.0800 0.3300 1.1550 0.8850 ;
        RECT 0.6750 0.2025 0.7950 0.3975 ;
        RECT 0.2775 0.6525 0.7800 0.7725 ;
        RECT 0.3750 0.2775 0.6750 0.3975 ;
        RECT 0.2550 0.2025 0.3750 0.3975 ;
    END
END DCCKN_0111


MACRO DCCKN_1100
    CLASS CORE ;
    FOREIGN DCCKN_1100 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.1400 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 1.9425 0.2775 2.1000 0.3975 ;
        RECT 1.9425 0.6525 2.1000 0.7725 ;
        RECT 1.6275 0.2775 1.9425 0.7725 ;
        RECT 1.4700 0.2775 1.6275 0.3975 ;
        RECT 1.4700 0.6525 1.6275 0.7725 ;
        VIA 1.9425 0.3375 VIA12_slot ;
        VIA 1.9425 0.7125 VIA12_slot ;
        VIA 1.6275 0.3375 VIA12_slot ;
        VIA 1.6275 0.7125 VIA12_slot ;
        END
    END ZN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1425 0.4725 3.4650 0.5475 ;
        RECT 0.0675 0.3675 0.1425 0.6825 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 6.4500 -0.0750 7.1400 0.0750 ;
        RECT 6.3525 -0.0750 6.4500 0.2625 ;
        RECT 3.5250 -0.0750 6.3525 0.0750 ;
        RECT 3.4050 -0.0750 3.5250 0.2925 ;
        RECT 3.1050 -0.0750 3.4050 0.0750 ;
        RECT 2.9850 -0.0750 3.1050 0.2025 ;
        RECT 2.6850 -0.0750 2.9850 0.0750 ;
        RECT 2.5650 -0.0750 2.6850 0.2025 ;
        RECT 2.2650 -0.0750 2.5650 0.0750 ;
        RECT 2.1450 -0.0750 2.2650 0.2025 ;
        RECT 1.8450 -0.0750 2.1450 0.0750 ;
        RECT 1.7250 -0.0750 1.8450 0.2025 ;
        RECT 1.4250 -0.0750 1.7250 0.0750 ;
        RECT 1.3050 -0.0750 1.4250 0.2025 ;
        RECT 1.0050 -0.0750 1.3050 0.0750 ;
        RECT 0.8850 -0.0750 1.0050 0.2025 ;
        RECT 0.5850 -0.0750 0.8850 0.0750 ;
        RECT 0.4650 -0.0750 0.5850 0.2025 ;
        RECT 0.1425 -0.0750 0.4650 0.0750 ;
        RECT 0.0675 -0.0750 0.1425 0.2475 ;
        RECT 0.0000 -0.0750 0.0675 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 7.0875 0.9750 7.1400 1.1250 ;
        RECT 6.9825 0.7725 7.0875 1.1250 ;
        RECT 6.8775 0.9750 6.9825 1.1250 ;
        RECT 6.7725 0.7725 6.8775 1.1250 ;
        RECT 6.6675 0.9750 6.7725 1.1250 ;
        RECT 6.5625 0.7725 6.6675 1.1250 ;
        RECT 6.4575 0.9750 6.5625 1.1250 ;
        RECT 6.3525 0.7725 6.4575 1.1250 ;
        RECT 6.2475 0.9750 6.3525 1.1250 ;
        RECT 6.1425 0.7725 6.2475 1.1250 ;
        RECT 6.0375 0.9750 6.1425 1.1250 ;
        RECT 5.9325 0.7725 6.0375 1.1250 ;
        RECT 5.8275 0.9750 5.9325 1.1250 ;
        RECT 5.7225 0.7725 5.8275 1.1250 ;
        RECT 5.6175 0.9750 5.7225 1.1250 ;
        RECT 5.5125 0.7725 5.6175 1.1250 ;
        RECT 5.4075 0.9750 5.5125 1.1250 ;
        RECT 5.3025 0.7725 5.4075 1.1250 ;
        RECT 5.1975 0.9750 5.3025 1.1250 ;
        RECT 5.0925 0.7725 5.1975 1.1250 ;
        RECT 4.9875 0.9750 5.0925 1.1250 ;
        RECT 4.8825 0.7725 4.9875 1.1250 ;
        RECT 4.7775 0.9750 4.8825 1.1250 ;
        RECT 4.6725 0.7725 4.7775 1.1250 ;
        RECT 4.5675 0.9750 4.6725 1.1250 ;
        RECT 4.4625 0.7725 4.5675 1.1250 ;
        RECT 4.3575 0.9750 4.4625 1.1250 ;
        RECT 4.2525 0.7725 4.3575 1.1250 ;
        RECT 4.1475 0.9750 4.2525 1.1250 ;
        RECT 4.0425 0.7725 4.1475 1.1250 ;
        RECT 3.9375 0.9750 4.0425 1.1250 ;
        RECT 3.8325 0.7725 3.9375 1.1250 ;
        RECT 3.5250 0.9750 3.8325 1.1250 ;
        RECT 3.4050 0.6600 3.5250 1.1250 ;
        RECT 3.1050 0.9750 3.4050 1.1250 ;
        RECT 2.9850 0.8475 3.1050 1.1250 ;
        RECT 2.6850 0.9750 2.9850 1.1250 ;
        RECT 2.5650 0.8475 2.6850 1.1250 ;
        RECT 2.2650 0.9750 2.5650 1.1250 ;
        RECT 2.1450 0.8475 2.2650 1.1250 ;
        RECT 1.8450 0.9750 2.1450 1.1250 ;
        RECT 1.7250 0.8475 1.8450 1.1250 ;
        RECT 1.4250 0.9750 1.7250 1.1250 ;
        RECT 1.3050 0.8475 1.4250 1.1250 ;
        RECT 1.0050 0.9750 1.3050 1.1250 ;
        RECT 0.8850 0.8475 1.0050 1.1250 ;
        RECT 0.5850 0.9750 0.8850 1.1250 ;
        RECT 0.4650 0.8475 0.5850 1.1250 ;
        RECT 0.1425 0.9750 0.4650 1.1250 ;
        RECT 0.0675 0.8025 0.1425 1.1250 ;
        RECT 0.0000 0.9750 0.0675 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 7.0050 0.8025 7.0650 0.8625 ;
        RECT 6.9000 0.6000 6.9600 0.6600 ;
        RECT 6.7950 0.8025 6.8550 0.8625 ;
        RECT 6.6900 0.6000 6.7500 0.6600 ;
        RECT 6.5850 0.1800 6.6450 0.2400 ;
        RECT 6.5850 0.8025 6.6450 0.8625 ;
        RECT 6.4800 0.3600 6.5400 0.4200 ;
        RECT 6.4800 0.6000 6.5400 0.6600 ;
        RECT 6.3750 0.1725 6.4350 0.2325 ;
        RECT 6.3750 0.8025 6.4350 0.8625 ;
        RECT 6.2700 0.5475 6.3300 0.6075 ;
        RECT 6.1650 0.8025 6.2250 0.8625 ;
        RECT 6.0600 0.5550 6.1200 0.6150 ;
        RECT 5.9550 0.8025 6.0150 0.8625 ;
        RECT 5.8500 0.5550 5.9100 0.6150 ;
        RECT 5.7450 0.8025 5.8050 0.8625 ;
        RECT 5.6400 0.5550 5.7000 0.6150 ;
        RECT 5.5350 0.8025 5.5950 0.8625 ;
        RECT 5.4300 0.5550 5.4900 0.6150 ;
        RECT 5.3250 0.8025 5.3850 0.8625 ;
        RECT 5.2200 0.5550 5.2800 0.6150 ;
        RECT 5.1150 0.8025 5.1750 0.8625 ;
        RECT 5.0100 0.5550 5.0700 0.6150 ;
        RECT 4.9050 0.8025 4.9650 0.8625 ;
        RECT 4.8000 0.5550 4.8600 0.6150 ;
        RECT 4.6950 0.8025 4.7550 0.8625 ;
        RECT 4.5900 0.5550 4.6500 0.6150 ;
        RECT 4.4850 0.8025 4.5450 0.8625 ;
        RECT 4.3800 0.5550 4.4400 0.6150 ;
        RECT 4.2750 0.8025 4.3350 0.8625 ;
        RECT 4.1700 0.5550 4.2300 0.6150 ;
        RECT 4.0650 0.8025 4.1250 0.8625 ;
        RECT 3.9600 0.5550 4.0200 0.6150 ;
        RECT 3.8550 0.8025 3.9150 0.8625 ;
        RECT 3.7500 0.5550 3.8100 0.6150 ;
        RECT 3.6450 0.7875 3.7050 0.8475 ;
        RECT 3.4350 0.2250 3.4950 0.2850 ;
        RECT 3.4350 0.6675 3.4950 0.7275 ;
        RECT 3.4350 0.8325 3.4950 0.8925 ;
        RECT 3.3300 0.4800 3.3900 0.5400 ;
        RECT 3.2250 0.3075 3.2850 0.3675 ;
        RECT 3.2250 0.6825 3.2850 0.7425 ;
        RECT 3.1200 0.4800 3.1800 0.5400 ;
        RECT 3.0150 0.1350 3.0750 0.1950 ;
        RECT 3.0150 0.8550 3.0750 0.9150 ;
        RECT 2.9100 0.4800 2.9700 0.5400 ;
        RECT 2.8050 0.3075 2.8650 0.3675 ;
        RECT 2.8050 0.6825 2.8650 0.7425 ;
        RECT 2.7000 0.4800 2.7600 0.5400 ;
        RECT 2.5950 0.1350 2.6550 0.1950 ;
        RECT 2.5950 0.8550 2.6550 0.9150 ;
        RECT 2.4900 0.4800 2.5500 0.5400 ;
        RECT 2.3850 0.3075 2.4450 0.3675 ;
        RECT 2.3850 0.6825 2.4450 0.7425 ;
        RECT 2.2800 0.4800 2.3400 0.5400 ;
        RECT 2.1750 0.1350 2.2350 0.1950 ;
        RECT 2.1750 0.8550 2.2350 0.9150 ;
        RECT 2.0700 0.4800 2.1300 0.5400 ;
        RECT 1.9650 0.3075 2.0250 0.3675 ;
        RECT 1.9650 0.6825 2.0250 0.7425 ;
        RECT 1.8600 0.4800 1.9200 0.5400 ;
        RECT 1.7550 0.1350 1.8150 0.1950 ;
        RECT 1.7550 0.8550 1.8150 0.9150 ;
        RECT 1.6500 0.4800 1.7100 0.5400 ;
        RECT 1.5450 0.3075 1.6050 0.3675 ;
        RECT 1.5450 0.6825 1.6050 0.7425 ;
        RECT 1.4400 0.4800 1.5000 0.5400 ;
        RECT 1.3350 0.1350 1.3950 0.1950 ;
        RECT 1.3350 0.8550 1.3950 0.9150 ;
        RECT 1.2300 0.4800 1.2900 0.5400 ;
        RECT 1.1250 0.3075 1.1850 0.3675 ;
        RECT 1.1250 0.6825 1.1850 0.7425 ;
        RECT 1.0200 0.4800 1.0800 0.5400 ;
        RECT 0.9150 0.1350 0.9750 0.1950 ;
        RECT 0.9150 0.8550 0.9750 0.9150 ;
        RECT 0.8100 0.4800 0.8700 0.5400 ;
        RECT 0.7050 0.3075 0.7650 0.3675 ;
        RECT 0.7050 0.6825 0.7650 0.7425 ;
        RECT 0.6000 0.4800 0.6600 0.5400 ;
        RECT 0.4950 0.1350 0.5550 0.1950 ;
        RECT 0.4950 0.8550 0.5550 0.9150 ;
        RECT 0.3900 0.4800 0.4500 0.5400 ;
        RECT 0.2850 0.3075 0.3450 0.3675 ;
        RECT 0.2850 0.6825 0.3450 0.7425 ;
        RECT 0.1800 0.4800 0.2400 0.5400 ;
        RECT 0.0750 0.1575 0.1350 0.2175 ;
        RECT 0.0750 0.8325 0.1350 0.8925 ;
        LAYER M1 ;
        RECT 6.7500 0.5850 7.0050 0.6675 ;
        RECT 6.6750 0.1725 6.7500 0.6675 ;
        RECT 6.5550 0.1725 6.6750 0.2475 ;
        RECT 6.3600 0.5775 6.6750 0.6675 ;
        RECT 3.6750 0.3525 6.5700 0.4275 ;
        RECT 6.2475 0.5400 6.3600 0.6675 ;
        RECT 3.8550 0.5400 6.2475 0.6150 ;
        RECT 3.7500 0.5250 3.8550 0.6450 ;
        RECT 3.6750 0.7575 3.7125 0.8850 ;
        RECT 3.6000 0.3525 3.6750 0.8850 ;
        RECT 0.2775 0.2775 3.3000 0.3975 ;
        RECT 0.2775 0.6525 3.3000 0.7725 ;
        LAYER M2 ;
        RECT 1.9725 0.2775 2.1000 0.3975 ;
        RECT 1.9725 0.6525 2.1000 0.7725 ;
        RECT 1.4700 0.2775 1.5975 0.3975 ;
        RECT 1.4700 0.6525 1.5975 0.7725 ;
    END
END DCCKN_1100


MACRO DEL025_1010
    CLASS CORE ;
    FOREIGN DEL025_1010 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.6300 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.5175 0.2175 0.5925 0.8325 ;
        RECT 0.4875 0.2175 0.5175 0.3825 ;
        RECT 0.4875 0.6675 0.5175 0.8325 ;
        END
    END Z
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.0375 0.4125 0.2400 0.6375 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.3750 -0.0750 0.6300 0.0750 ;
        RECT 0.2550 -0.0750 0.3750 0.1875 ;
        RECT 0.0000 -0.0750 0.2550 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.3750 0.9750 0.6300 1.1250 ;
        RECT 0.2550 0.8625 0.3750 1.1250 ;
        RECT 0.0000 0.9750 0.2550 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 0.4950 0.2700 0.5550 0.3300 ;
        RECT 0.4950 0.7200 0.5550 0.7800 ;
        RECT 0.3825 0.4800 0.4425 0.5400 ;
        RECT 0.2850 0.1275 0.3450 0.1875 ;
        RECT 0.2850 0.8625 0.3450 0.9225 ;
        RECT 0.1800 0.4875 0.2400 0.5475 ;
        RECT 0.0750 0.1725 0.1350 0.2325 ;
        RECT 0.0750 0.8025 0.1350 0.8625 ;
        LAYER M1 ;
        RECT 0.3900 0.4500 0.4425 0.5700 ;
        RECT 0.3150 0.2625 0.3900 0.7875 ;
        RECT 0.1575 0.2625 0.3150 0.3375 ;
        RECT 0.1575 0.7125 0.3150 0.7875 ;
        RECT 0.0525 0.1500 0.1575 0.3375 ;
        RECT 0.0525 0.7125 0.1575 0.8850 ;
    END
END DEL025_1010


MACRO DEL150M_1010
    CLASS CORE ;
    FOREIGN DEL150M_1010 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.4100 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 4.2975 0.2175 4.3725 0.8325 ;
        RECT 4.2675 0.2175 4.2975 0.3825 ;
        RECT 4.2675 0.6675 4.2975 0.8325 ;
        END
    END Z
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.0375 0.4050 0.2400 0.6375 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 4.1550 -0.0750 4.4100 0.0750 ;
        RECT 4.0350 -0.0750 4.1550 0.1800 ;
        RECT 2.6850 -0.0750 4.0350 0.0750 ;
        RECT 2.5650 -0.0750 2.6850 0.2400 ;
        RECT 0.3750 -0.0750 2.5650 0.0750 ;
        RECT 0.2550 -0.0750 0.3750 0.1800 ;
        RECT 0.0000 -0.0750 0.2550 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 4.1550 0.9750 4.4100 1.1250 ;
        RECT 4.0350 0.8625 4.1550 1.1250 ;
        RECT 2.6850 0.9750 4.0350 1.1250 ;
        RECT 2.5650 0.7950 2.6850 1.1250 ;
        RECT 0.3750 0.9750 2.5650 1.1250 ;
        RECT 0.2550 0.8625 0.3750 1.1250 ;
        RECT 0.0000 0.9750 0.2550 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 4.2750 0.2775 4.3350 0.3375 ;
        RECT 4.2750 0.7275 4.3350 0.7875 ;
        RECT 4.1625 0.4950 4.2225 0.5550 ;
        RECT 4.0650 0.1200 4.1250 0.1800 ;
        RECT 4.0650 0.8625 4.1250 0.9225 ;
        RECT 3.9525 0.4725 4.0125 0.5325 ;
        RECT 3.8550 0.2175 3.9150 0.2775 ;
        RECT 3.8550 0.7950 3.9150 0.8550 ;
        RECT 3.6450 0.2175 3.7050 0.2775 ;
        RECT 3.6450 0.7950 3.7050 0.8550 ;
        RECT 3.5475 0.4725 3.6075 0.5325 ;
        RECT 3.4350 0.2325 3.4950 0.2925 ;
        RECT 3.4350 0.7800 3.4950 0.8400 ;
        RECT 3.2250 0.1950 3.2850 0.2550 ;
        RECT 3.2250 0.7425 3.2850 0.8025 ;
        RECT 3.1125 0.4650 3.1725 0.5250 ;
        RECT 3.0150 0.1875 3.0750 0.2475 ;
        RECT 3.0150 0.7425 3.0750 0.8025 ;
        RECT 2.8050 0.1875 2.8650 0.2475 ;
        RECT 2.8050 0.7425 2.8650 0.8025 ;
        RECT 2.7000 0.4650 2.7600 0.5250 ;
        RECT 2.5950 0.1800 2.6550 0.2400 ;
        RECT 2.5950 0.7950 2.6550 0.8550 ;
        RECT 2.4900 0.4950 2.5500 0.5550 ;
        RECT 2.3850 0.2550 2.4450 0.3150 ;
        RECT 2.3850 0.7575 2.4450 0.8175 ;
        RECT 2.1750 0.2475 2.2350 0.3075 ;
        RECT 2.1750 0.7725 2.2350 0.8325 ;
        RECT 2.0775 0.4875 2.1375 0.5475 ;
        RECT 1.9650 0.1950 2.0250 0.2550 ;
        RECT 1.9650 0.7875 2.0250 0.8475 ;
        RECT 1.7550 0.1950 1.8150 0.2550 ;
        RECT 1.7550 0.7875 1.8150 0.8475 ;
        RECT 1.6575 0.4875 1.7175 0.5475 ;
        RECT 1.5450 0.2325 1.6050 0.2925 ;
        RECT 1.5450 0.7800 1.6050 0.8400 ;
        RECT 1.3350 0.1875 1.3950 0.2475 ;
        RECT 1.3350 0.7800 1.3950 0.8400 ;
        RECT 1.2225 0.4875 1.2825 0.5475 ;
        RECT 1.1250 0.1875 1.1850 0.2475 ;
        RECT 1.1250 0.7725 1.1850 0.8325 ;
        RECT 0.9150 0.1875 0.9750 0.2475 ;
        RECT 0.9150 0.7725 0.9750 0.8325 ;
        RECT 0.8025 0.4875 0.8625 0.5475 ;
        RECT 0.7050 0.2100 0.7650 0.2700 ;
        RECT 0.7050 0.7725 0.7650 0.8325 ;
        RECT 0.4950 0.2100 0.5550 0.2700 ;
        RECT 0.4950 0.7575 0.5550 0.8175 ;
        RECT 0.3900 0.4650 0.4500 0.5250 ;
        RECT 0.2850 0.1200 0.3450 0.1800 ;
        RECT 0.2850 0.8625 0.3450 0.9225 ;
        RECT 0.1800 0.4650 0.2400 0.5250 ;
        RECT 0.0750 0.1725 0.1350 0.2325 ;
        RECT 0.0750 0.7500 0.1350 0.8100 ;
        LAYER M1 ;
        RECT 4.1925 0.4650 4.2225 0.6075 ;
        RECT 4.0875 0.2850 4.1925 0.6075 ;
        RECT 3.8925 0.4350 4.0125 0.6975 ;
        RECT 3.8175 0.1875 3.9450 0.2925 ;
        RECT 3.8175 0.7800 3.9450 0.8925 ;
        RECT 3.7425 0.1875 3.8175 0.8925 ;
        RECT 3.6150 0.1875 3.7425 0.3000 ;
        RECT 3.6150 0.7800 3.7425 0.8925 ;
        RECT 3.5475 0.4275 3.6675 0.6900 ;
        RECT 3.4725 0.2025 3.4950 0.3300 ;
        RECT 3.4725 0.7500 3.4950 0.8700 ;
        RECT 3.3975 0.2025 3.4725 0.8700 ;
        RECT 3.2475 0.1725 3.3225 0.8325 ;
        RECT 3.1950 0.1725 3.2475 0.2775 ;
        RECT 3.2250 0.7125 3.2475 0.8325 ;
        RECT 3.0525 0.3600 3.1725 0.6225 ;
        RECT 2.9775 0.1650 3.1050 0.2700 ;
        RECT 2.9775 0.7200 3.1050 0.8250 ;
        RECT 2.9025 0.1650 2.9775 0.8250 ;
        RECT 2.7750 0.1650 2.9025 0.2775 ;
        RECT 2.7750 0.7200 2.9025 0.8250 ;
        RECT 2.6775 0.3600 2.8275 0.5925 ;
        RECT 2.4225 0.4425 2.5725 0.6525 ;
        RECT 2.3475 0.2175 2.4525 0.3450 ;
        RECT 2.3475 0.7275 2.4525 0.8625 ;
        RECT 2.2725 0.2175 2.3475 0.8625 ;
        RECT 2.1450 0.2175 2.2725 0.3300 ;
        RECT 2.1450 0.7575 2.2725 0.8625 ;
        RECT 2.0775 0.4125 2.1975 0.6750 ;
        RECT 1.9275 0.1800 2.0550 0.2850 ;
        RECT 1.9275 0.7575 2.0550 0.8700 ;
        RECT 1.8525 0.1800 1.9275 0.8700 ;
        RECT 1.7250 0.1800 1.8525 0.2925 ;
        RECT 1.7250 0.7575 1.8525 0.8700 ;
        RECT 1.6575 0.4125 1.7775 0.6750 ;
        RECT 1.5825 0.2025 1.6050 0.3300 ;
        RECT 1.5825 0.7500 1.6050 0.8700 ;
        RECT 1.5075 0.2025 1.5825 0.8700 ;
        RECT 1.3575 0.1800 1.4325 0.8700 ;
        RECT 1.3050 0.1800 1.3575 0.2850 ;
        RECT 1.3350 0.7275 1.3575 0.8700 ;
        RECT 1.1625 0.3600 1.2825 0.6225 ;
        RECT 1.0800 0.1650 1.2075 0.2700 ;
        RECT 1.0800 0.7425 1.2075 0.8550 ;
        RECT 1.0050 0.1650 1.0800 0.8550 ;
        RECT 0.8775 0.1650 1.0050 0.2775 ;
        RECT 0.8775 0.7425 1.0050 0.8550 ;
        RECT 0.7425 0.3600 0.8625 0.6225 ;
        RECT 0.6675 0.1800 0.7950 0.2850 ;
        RECT 0.6675 0.7575 0.7950 0.8625 ;
        RECT 0.5925 0.1800 0.6675 0.8625 ;
        RECT 0.4875 0.1800 0.5925 0.3000 ;
        RECT 0.4875 0.7275 0.5925 0.8625 ;
        RECT 0.3900 0.3750 0.5175 0.5400 ;
        RECT 0.3150 0.2550 0.3900 0.7875 ;
        RECT 0.1575 0.2550 0.3150 0.3300 ;
        RECT 0.1575 0.7125 0.3150 0.7875 ;
        RECT 0.0525 0.1500 0.1575 0.3300 ;
        RECT 0.0525 0.7125 0.1575 0.8550 ;
        LAYER VIA1 ;
        RECT 4.1025 0.4125 4.1775 0.4875 ;
        RECT 3.9150 0.5625 3.9900 0.6375 ;
        RECT 3.5775 0.5625 3.6525 0.6375 ;
        RECT 3.3975 0.4125 3.4725 0.4875 ;
        RECT 3.2475 0.5625 3.3225 0.6375 ;
        RECT 3.0675 0.4125 3.1425 0.4875 ;
        RECT 2.7150 0.4125 2.7900 0.4875 ;
        RECT 2.4600 0.5625 2.5350 0.6375 ;
        RECT 2.0925 0.5625 2.1675 0.6375 ;
        RECT 1.6800 0.5625 1.7550 0.6375 ;
        RECT 1.5075 0.4125 1.5825 0.4875 ;
        RECT 1.3575 0.5625 1.4325 0.6375 ;
        RECT 1.1775 0.4125 1.2525 0.4875 ;
        RECT 0.7725 0.4125 0.8475 0.4875 ;
        RECT 0.4050 0.4125 0.4800 0.4875 ;
        LAYER M2 ;
        RECT 3.3525 0.4125 4.2450 0.4875 ;
        RECT 3.1875 0.5625 4.0350 0.6375 ;
        RECT 1.4400 0.4125 3.1875 0.4875 ;
        RECT 1.3125 0.5625 2.5800 0.6375 ;
        RECT 0.3600 0.4125 1.3050 0.4875 ;
    END
END DEL150M_1010


MACRO DFCNQ_0011
    CLASS CORE ;
    FOREIGN DFCNQ_0011 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.2000 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 4.0875 0.3150 4.1625 0.7350 ;
        RECT 3.9225 0.3150 4.0875 0.3900 ;
        RECT 3.9225 0.6600 4.0875 0.7350 ;
        RECT 3.8475 0.2175 3.9225 0.3900 ;
        RECT 3.8475 0.6600 3.9225 0.8325 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.4500 0.5625 0.9150 0.6375 ;
        VIA 0.7125 0.6000 VIA12_square ;
        END
    END D
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.0675 0.4125 0.6225 0.4875 ;
        VIA 0.1800 0.4500 VIA12_square ;
        END
    END CP
    PIN CDN
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 3.4575 0.1125 3.5325 0.5775 ;
        RECT 1.7550 0.1125 3.4575 0.1875 ;
        RECT 1.6500 0.1125 1.7550 0.5250 ;
        VIA 3.4950 0.4950 VIA12_square ;
        VIA 1.7025 0.4425 VIA12_square ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 4.1550 -0.0750 4.2000 0.0750 ;
        RECT 4.0350 -0.0750 4.1550 0.2400 ;
        RECT 3.7350 -0.0750 4.0350 0.0750 ;
        RECT 3.6150 -0.0750 3.7350 0.1800 ;
        RECT 3.1050 -0.0750 3.6150 0.0750 ;
        RECT 2.9850 -0.0750 3.1050 0.2175 ;
        RECT 2.0550 -0.0750 2.9850 0.0750 ;
        RECT 1.9350 -0.0750 2.0550 0.1800 ;
        RECT 0.7875 -0.0750 1.9350 0.0750 ;
        RECT 0.6825 -0.0750 0.7875 0.2400 ;
        RECT 0.3750 -0.0750 0.6825 0.0750 ;
        RECT 0.2550 -0.0750 0.3750 0.1875 ;
        RECT 0.0000 -0.0750 0.2550 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 4.1475 0.9750 4.2000 1.1250 ;
        RECT 4.0425 0.8100 4.1475 1.1250 ;
        RECT 3.7350 0.9750 4.0425 1.1250 ;
        RECT 3.6150 0.8475 3.7350 1.1250 ;
        RECT 3.3000 0.9750 3.6150 1.1250 ;
        RECT 3.2250 0.8325 3.3000 1.1250 ;
        RECT 2.0550 0.9750 3.2250 1.1250 ;
        RECT 1.9500 0.8100 2.0550 1.1250 ;
        RECT 1.6350 0.9750 1.9500 1.1250 ;
        RECT 1.5150 0.8325 1.6350 1.1250 ;
        RECT 0.7725 0.9750 1.5150 1.1250 ;
        RECT 0.6975 0.7950 0.7725 1.1250 ;
        RECT 0.3750 0.9750 0.6975 1.1250 ;
        RECT 0.2550 0.8625 0.3750 1.1250 ;
        RECT 0.0000 0.9750 0.2550 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 4.0650 0.1575 4.1250 0.2175 ;
        RECT 4.0650 0.8325 4.1250 0.8925 ;
        RECT 3.9525 0.4950 4.0125 0.5550 ;
        RECT 3.8550 0.2700 3.9150 0.3300 ;
        RECT 3.8550 0.7200 3.9150 0.7800 ;
        RECT 3.7500 0.4950 3.8100 0.5550 ;
        RECT 3.6450 0.1200 3.7050 0.1800 ;
        RECT 3.6450 0.8700 3.7050 0.9300 ;
        RECT 3.5400 0.4725 3.6000 0.5325 ;
        RECT 3.4350 0.8325 3.4950 0.8925 ;
        RECT 3.3225 0.4950 3.3825 0.5550 ;
        RECT 3.2250 0.2850 3.2850 0.3450 ;
        RECT 3.2250 0.8625 3.2850 0.9225 ;
        RECT 3.1200 0.4875 3.1800 0.5475 ;
        RECT 3.0150 0.1575 3.0750 0.2175 ;
        RECT 3.0150 0.8325 3.0750 0.8925 ;
        RECT 2.9100 0.4875 2.9700 0.5475 ;
        RECT 2.7000 0.5250 2.7600 0.5850 ;
        RECT 2.5950 0.1725 2.6550 0.2325 ;
        RECT 2.5950 0.8325 2.6550 0.8925 ;
        RECT 2.4900 0.3750 2.5500 0.4350 ;
        RECT 2.3850 0.1725 2.4450 0.2325 ;
        RECT 2.3850 0.7350 2.4450 0.7950 ;
        RECT 2.2800 0.5175 2.3400 0.5775 ;
        RECT 2.1750 0.1575 2.2350 0.2175 ;
        RECT 2.1750 0.8175 2.2350 0.8775 ;
        RECT 2.0700 0.3750 2.1300 0.4350 ;
        RECT 1.9650 0.1200 2.0250 0.1800 ;
        RECT 1.9650 0.8400 2.0250 0.9000 ;
        RECT 1.8600 0.5400 1.9200 0.6000 ;
        RECT 1.7550 0.8325 1.8150 0.8925 ;
        RECT 1.6500 0.4800 1.7100 0.5400 ;
        RECT 1.5450 0.8325 1.6050 0.8925 ;
        RECT 1.4400 0.4575 1.5000 0.5175 ;
        RECT 1.3350 0.1800 1.3950 0.2400 ;
        RECT 1.3350 0.8100 1.3950 0.8700 ;
        RECT 1.2300 0.5025 1.2900 0.5625 ;
        RECT 1.1250 0.1725 1.1850 0.2325 ;
        RECT 1.1250 0.8025 1.1850 0.8625 ;
        RECT 1.0200 0.3600 1.0800 0.4200 ;
        RECT 0.9150 0.1725 0.9750 0.2325 ;
        RECT 0.8100 0.5250 0.8700 0.5850 ;
        RECT 0.7050 0.1575 0.7650 0.2175 ;
        RECT 0.7050 0.8325 0.7650 0.8925 ;
        RECT 0.4950 0.2775 0.5550 0.3375 ;
        RECT 0.4950 0.7350 0.5550 0.7950 ;
        RECT 0.3900 0.4650 0.4500 0.5250 ;
        RECT 0.2850 0.1200 0.3450 0.1800 ;
        RECT 0.2850 0.8700 0.3450 0.9300 ;
        RECT 0.1800 0.4875 0.2400 0.5475 ;
        RECT 0.0750 0.2400 0.1350 0.3000 ;
        RECT 0.0750 0.7500 0.1350 0.8100 ;
        LAYER M1 ;
        RECT 3.7575 0.4650 4.0125 0.5850 ;
        RECT 3.6825 0.2625 3.7575 0.7725 ;
        RECT 3.3600 0.2625 3.6825 0.3375 ;
        RECT 3.5400 0.6975 3.6825 0.7725 ;
        RECT 3.4575 0.4125 3.6075 0.6225 ;
        RECT 3.4650 0.6975 3.5400 0.9000 ;
        RECT 3.4050 0.8100 3.4650 0.9000 ;
        RECT 3.3075 0.4650 3.3825 0.7275 ;
        RECT 3.2850 0.2625 3.3600 0.3525 ;
        RECT 3.1125 0.6525 3.3075 0.7275 ;
        RECT 3.2325 0.2775 3.2850 0.3525 ;
        RECT 3.1575 0.2775 3.2325 0.5775 ;
        RECT 2.9100 0.4575 3.1575 0.5775 ;
        RECT 2.5500 0.8250 3.1200 0.9000 ;
        RECT 3.0375 0.6525 3.1125 0.7500 ;
        RECT 2.4450 0.6750 3.0375 0.7500 ;
        RECT 2.8800 0.2925 2.9700 0.3825 ;
        RECT 2.7900 0.1500 2.8800 0.3825 ;
        RECT 2.5725 0.1500 2.7900 0.2550 ;
        RECT 2.2500 0.5175 2.7900 0.5925 ;
        RECT 2.4150 0.3300 2.7150 0.4350 ;
        RECT 2.3400 0.1500 2.4675 0.2550 ;
        RECT 2.3700 0.6750 2.4450 0.8400 ;
        RECT 2.2350 0.1500 2.3400 0.4425 ;
        RECT 2.2125 0.8100 2.2650 0.8850 ;
        RECT 2.1450 0.1500 2.2350 0.2550 ;
        RECT 2.1375 0.6600 2.2125 0.8850 ;
        RECT 2.0475 0.3300 2.1600 0.4350 ;
        RECT 2.0250 0.6600 2.1375 0.7350 ;
        RECT 1.9725 0.2550 2.0475 0.4350 ;
        RECT 1.8600 0.5100 2.0250 0.7350 ;
        RECT 1.8450 0.2550 1.9725 0.3300 ;
        RECT 1.7700 0.1950 1.8450 0.3300 ;
        RECT 1.7850 0.8175 1.8450 0.9000 ;
        RECT 1.6200 0.4050 1.7850 0.6000 ;
        RECT 1.7100 0.6825 1.7850 0.9000 ;
        RECT 1.4850 0.1950 1.7700 0.2700 ;
        RECT 1.4400 0.6825 1.7100 0.7575 ;
        RECT 1.4250 0.3450 1.5300 0.6075 ;
        RECT 1.3350 0.1500 1.4850 0.2700 ;
        RECT 1.3350 0.6825 1.4400 0.9000 ;
        RECT 0.6000 0.3450 1.4250 0.4200 ;
        RECT 1.0200 0.4950 1.3200 0.5700 ;
        RECT 1.0950 0.6450 1.2600 0.9000 ;
        RECT 0.8925 0.1500 1.2300 0.2550 ;
        RECT 0.9450 0.4950 1.0200 0.9000 ;
        RECT 0.8550 0.7800 0.9450 0.9000 ;
        RECT 0.6750 0.4950 0.8700 0.6900 ;
        RECT 0.5625 0.2475 0.6000 0.7200 ;
        RECT 0.5250 0.2475 0.5625 0.8400 ;
        RECT 0.4875 0.2475 0.5250 0.3675 ;
        RECT 0.4875 0.6450 0.5250 0.8400 ;
        RECT 0.4125 0.4350 0.4500 0.5550 ;
        RECT 0.3375 0.2625 0.4125 0.7875 ;
        RECT 0.1425 0.2625 0.3375 0.3375 ;
        RECT 0.1425 0.7125 0.3375 0.7875 ;
        RECT 0.0975 0.4125 0.2625 0.6375 ;
        RECT 0.0675 0.2025 0.1425 0.3375 ;
        RECT 0.0675 0.7125 0.1425 0.8475 ;
        LAYER VIA1 ;
        RECT 2.8500 0.3000 2.9250 0.3750 ;
        RECT 2.8050 0.6750 2.8800 0.7500 ;
        RECT 2.6550 0.5175 2.7300 0.5925 ;
        RECT 2.4675 0.3450 2.5425 0.4200 ;
        RECT 2.2500 0.3300 2.3250 0.4050 ;
        RECT 1.9050 0.5100 1.9800 0.5850 ;
        RECT 1.4325 0.4875 1.5075 0.5625 ;
        RECT 1.3800 0.1950 1.4550 0.2700 ;
        RECT 1.1400 0.6600 1.2150 0.7350 ;
        RECT 0.9000 0.8025 0.9750 0.8775 ;
        RECT 0.2925 0.7125 0.3675 0.7875 ;
        LAYER M2 ;
        RECT 2.8800 0.2925 2.9700 0.3975 ;
        RECT 2.8050 0.2925 2.8800 0.7950 ;
        RECT 2.6550 0.4725 2.7300 0.8850 ;
        RECT 1.0200 0.8100 2.6550 0.8850 ;
        RECT 2.5125 0.3150 2.5800 0.4500 ;
        RECT 2.4375 0.3150 2.5125 0.7350 ;
        RECT 1.5075 0.6600 2.4375 0.7350 ;
        RECT 2.2125 0.3150 2.3625 0.4200 ;
        RECT 2.1375 0.3150 2.2125 0.5850 ;
        RECT 1.9650 0.5100 2.1375 0.5850 ;
        RECT 1.8600 0.4800 1.9650 0.5850 ;
        RECT 1.4325 0.4425 1.5075 0.7350 ;
        RECT 1.2600 0.1950 1.5000 0.2700 ;
        RECT 1.1850 0.1950 1.2600 0.7350 ;
        RECT 1.0950 0.6600 1.1850 0.7350 ;
        RECT 0.8550 0.7950 1.0200 0.8850 ;
        RECT 0.4650 0.7950 0.8550 0.8700 ;
        RECT 0.3900 0.7125 0.4650 0.8700 ;
        RECT 0.2475 0.7125 0.3900 0.7875 ;
    END
END DFCNQ_0011


MACRO DFCNQ_0111
    CLASS CORE ;
    FOREIGN DFCNQ_0111 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.8300 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 4.1475 0.2325 4.4625 0.7350 ;
        VIA 4.3050 0.3150 VIA12_slot ;
        VIA 4.3050 0.6525 VIA12_slot ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.4500 0.5625 0.9150 0.6375 ;
        VIA 0.7125 0.6000 VIA12_square ;
        END
    END D
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.0675 0.4125 0.6225 0.4875 ;
        VIA 0.1800 0.4500 VIA12_square ;
        END
    END CP
    PIN CDN
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 3.7275 0.1125 3.8025 0.7875 ;
        RECT 1.7550 0.1125 3.7275 0.1875 ;
        RECT 3.2550 0.7125 3.7275 0.7875 ;
        RECT 3.1800 0.4725 3.2550 0.7875 ;
        RECT 1.6800 0.1125 1.7550 0.4275 ;
        RECT 1.5825 0.3225 1.6800 0.4275 ;
        VIA 3.7650 0.5325 VIA12_square ;
        VIA 3.2175 0.5625 VIA12_square ;
        VIA 1.6725 0.3750 VIA12_square ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 4.7700 -0.0750 4.8300 0.0750 ;
        RECT 4.6950 -0.0750 4.7700 0.2850 ;
        RECT 4.3650 -0.0750 4.6950 0.0750 ;
        RECT 4.2450 -0.0750 4.3650 0.1875 ;
        RECT 3.9450 -0.0750 4.2450 0.0750 ;
        RECT 3.8400 -0.0750 3.9450 0.2250 ;
        RECT 3.0900 -0.0750 3.8400 0.0750 ;
        RECT 3.0000 -0.0750 3.0900 0.2475 ;
        RECT 2.0400 -0.0750 3.0000 0.0750 ;
        RECT 1.9650 -0.0750 2.0400 0.2550 ;
        RECT 0.7875 -0.0750 1.9650 0.0750 ;
        RECT 0.6825 -0.0750 0.7875 0.2400 ;
        RECT 0.3750 -0.0750 0.6825 0.0750 ;
        RECT 0.2550 -0.0750 0.3750 0.1875 ;
        RECT 0.0000 -0.0750 0.2550 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 4.7625 0.9750 4.8300 1.1250 ;
        RECT 4.6875 0.7500 4.7625 1.1250 ;
        RECT 4.3650 0.9750 4.6875 1.1250 ;
        RECT 4.2450 0.8175 4.3650 1.1250 ;
        RECT 3.9450 0.9750 4.2450 1.1250 ;
        RECT 3.8250 0.8700 3.9450 1.1250 ;
        RECT 3.5250 0.9750 3.8250 1.1250 ;
        RECT 3.4050 0.8700 3.5250 1.1250 ;
        RECT 3.1050 0.9750 3.4050 1.1250 ;
        RECT 2.9850 0.8700 3.1050 1.1250 ;
        RECT 2.0250 0.9750 2.9850 1.1250 ;
        RECT 1.9500 0.8400 2.0250 1.1250 ;
        RECT 1.6050 0.9750 1.9500 1.1250 ;
        RECT 1.5300 0.8025 1.6050 1.1250 ;
        RECT 0.7725 0.9750 1.5300 1.1250 ;
        RECT 0.6975 0.7950 0.7725 1.1250 ;
        RECT 0.3750 0.9750 0.6975 1.1250 ;
        RECT 0.2550 0.8625 0.3750 1.1250 ;
        RECT 0.0000 0.9750 0.2550 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 4.6950 0.1950 4.7550 0.2550 ;
        RECT 4.6950 0.7950 4.7550 0.8550 ;
        RECT 4.5900 0.4725 4.6500 0.5325 ;
        RECT 4.4850 0.2850 4.5450 0.3450 ;
        RECT 4.4850 0.6525 4.5450 0.7125 ;
        RECT 4.3800 0.4725 4.4400 0.5325 ;
        RECT 4.2750 0.1275 4.3350 0.1875 ;
        RECT 4.2750 0.8325 4.3350 0.8925 ;
        RECT 4.1700 0.4725 4.2300 0.5325 ;
        RECT 4.0650 0.2700 4.1250 0.3300 ;
        RECT 4.0650 0.6525 4.1250 0.7125 ;
        RECT 3.9600 0.4725 4.0200 0.5325 ;
        RECT 3.8550 0.1350 3.9150 0.1950 ;
        RECT 3.8550 0.8700 3.9150 0.9300 ;
        RECT 3.7500 0.4950 3.8100 0.5550 ;
        RECT 3.6450 0.1575 3.7050 0.2175 ;
        RECT 3.6450 0.7275 3.7050 0.7875 ;
        RECT 3.5400 0.4875 3.6000 0.5475 ;
        RECT 3.4350 0.3075 3.4950 0.3675 ;
        RECT 3.4350 0.8700 3.4950 0.9300 ;
        RECT 3.3375 0.4875 3.3975 0.5475 ;
        RECT 3.2250 0.1575 3.2850 0.2175 ;
        RECT 3.2250 0.7275 3.2850 0.7875 ;
        RECT 3.1200 0.4875 3.1800 0.5475 ;
        RECT 3.0150 0.1575 3.0750 0.2175 ;
        RECT 3.0150 0.8700 3.0750 0.9300 ;
        RECT 2.9100 0.4800 2.9700 0.5400 ;
        RECT 2.8050 0.8175 2.8650 0.8775 ;
        RECT 2.7000 0.4800 2.7600 0.5400 ;
        RECT 2.5950 0.1725 2.6550 0.2325 ;
        RECT 2.5950 0.8100 2.6550 0.8700 ;
        RECT 2.4900 0.4200 2.5500 0.4800 ;
        RECT 2.3850 0.1800 2.4450 0.2400 ;
        RECT 2.3850 0.8100 2.4450 0.8700 ;
        RECT 2.2875 0.5625 2.3475 0.6225 ;
        RECT 2.1750 0.1800 2.2350 0.2400 ;
        RECT 2.1750 0.8100 2.2350 0.8700 ;
        RECT 2.0625 0.4200 2.1225 0.4800 ;
        RECT 1.9650 0.1650 2.0250 0.2250 ;
        RECT 1.9650 0.8700 2.0250 0.9300 ;
        RECT 1.8600 0.5625 1.9200 0.6225 ;
        RECT 1.7550 0.8325 1.8150 0.8925 ;
        RECT 1.6500 0.4500 1.7100 0.5100 ;
        RECT 1.5450 0.8325 1.6050 0.8925 ;
        RECT 1.4400 0.4350 1.5000 0.4950 ;
        RECT 1.3350 0.1800 1.3950 0.2400 ;
        RECT 1.3350 0.8100 1.3950 0.8700 ;
        RECT 1.2225 0.5025 1.2825 0.5625 ;
        RECT 1.1250 0.1725 1.1850 0.2325 ;
        RECT 1.1250 0.8025 1.1850 0.8625 ;
        RECT 1.0200 0.3525 1.0800 0.4125 ;
        RECT 0.9150 0.1725 0.9750 0.2325 ;
        RECT 0.8100 0.5250 0.8700 0.5850 ;
        RECT 0.7050 0.1575 0.7650 0.2175 ;
        RECT 0.7050 0.8325 0.7650 0.8925 ;
        RECT 0.4950 0.2775 0.5550 0.3375 ;
        RECT 0.4950 0.7350 0.5550 0.7950 ;
        RECT 0.3900 0.4650 0.4500 0.5250 ;
        RECT 0.2850 0.1200 0.3450 0.1800 ;
        RECT 0.2850 0.8700 0.3450 0.9300 ;
        RECT 0.1800 0.4875 0.2400 0.5475 ;
        RECT 0.0750 0.2400 0.1350 0.3000 ;
        RECT 0.0750 0.7500 0.1350 0.8100 ;
        LAYER M1 ;
        RECT 4.5600 0.4350 4.6800 0.5400 ;
        RECT 4.1475 0.2625 4.5750 0.3600 ;
        RECT 4.0650 0.6150 4.5675 0.7425 ;
        RECT 3.9900 0.4650 4.5600 0.5400 ;
        RECT 4.0650 0.2400 4.1475 0.3600 ;
        RECT 3.9150 0.3000 3.9900 0.7950 ;
        RECT 3.3900 0.3000 3.9150 0.3750 ;
        RECT 3.0450 0.7200 3.9150 0.7950 ;
        RECT 3.6750 0.4500 3.8400 0.6450 ;
        RECT 3.1950 0.1500 3.7350 0.2250 ;
        RECT 3.3375 0.4500 3.6000 0.5775 ;
        RECT 3.1200 0.3675 3.2625 0.6450 ;
        RECT 2.9700 0.4575 3.0450 0.7950 ;
        RECT 2.8800 0.4575 2.9700 0.5625 ;
        RECT 2.5950 0.7800 2.8950 0.9000 ;
        RECT 2.6775 0.4575 2.7825 0.6750 ;
        RECT 2.6550 0.1500 2.7600 0.3825 ;
        RECT 2.2575 0.5625 2.6775 0.6750 ;
        RECT 2.5200 0.1500 2.6550 0.2850 ;
        RECT 2.3550 0.3600 2.5800 0.4875 ;
        RECT 2.3100 0.7500 2.5200 0.9000 ;
        RECT 2.2800 0.1500 2.4450 0.2700 ;
        RECT 2.2575 0.4125 2.3550 0.4875 ;
        RECT 2.1150 0.1500 2.2800 0.3375 ;
        RECT 2.1750 0.7800 2.2350 0.9000 ;
        RECT 2.1000 0.6600 2.1750 0.9000 ;
        RECT 1.8900 0.4125 2.1525 0.4875 ;
        RECT 1.9950 0.6600 2.1000 0.7350 ;
        RECT 1.8300 0.5625 1.9950 0.7350 ;
        RECT 1.8150 0.1500 1.8900 0.4875 ;
        RECT 1.7550 0.8175 1.8450 0.9000 ;
        RECT 1.4700 0.1500 1.8150 0.2250 ;
        RECT 1.6800 0.6225 1.7550 0.9000 ;
        RECT 1.5975 0.3000 1.7400 0.5475 ;
        RECT 1.4550 0.6225 1.6800 0.6975 ;
        RECT 1.4175 0.3450 1.5225 0.5475 ;
        RECT 1.3050 0.1500 1.4700 0.2700 ;
        RECT 1.3800 0.6225 1.4550 0.9000 ;
        RECT 0.6000 0.3450 1.4175 0.4200 ;
        RECT 1.3350 0.7575 1.3800 0.9000 ;
        RECT 1.0200 0.4950 1.3125 0.5700 ;
        RECT 1.0950 0.6450 1.2600 0.9000 ;
        RECT 0.8925 0.1500 1.2300 0.2550 ;
        RECT 0.9450 0.4950 1.0200 0.9000 ;
        RECT 0.8550 0.7800 0.9450 0.9000 ;
        RECT 0.6750 0.4950 0.8700 0.6900 ;
        RECT 0.5625 0.2475 0.6000 0.7200 ;
        RECT 0.5250 0.2475 0.5625 0.8400 ;
        RECT 0.4875 0.2475 0.5250 0.3675 ;
        RECT 0.4875 0.6450 0.5250 0.8400 ;
        RECT 0.4125 0.4350 0.4500 0.5550 ;
        RECT 0.3375 0.2625 0.4125 0.7875 ;
        RECT 0.1425 0.2625 0.3375 0.3375 ;
        RECT 0.1425 0.7125 0.3375 0.7875 ;
        RECT 0.0975 0.4125 0.2625 0.6375 ;
        RECT 0.0675 0.2025 0.1425 0.3375 ;
        RECT 0.0675 0.7125 0.1425 0.8475 ;
        LAYER VIA1 ;
        RECT 3.4275 0.4725 3.5025 0.5475 ;
        RECT 2.6700 0.2625 2.7450 0.3375 ;
        RECT 2.4300 0.3975 2.5050 0.4725 ;
        RECT 2.4075 0.7950 2.4825 0.8700 ;
        RECT 2.3175 0.6000 2.3925 0.6750 ;
        RECT 2.1600 0.2625 2.2350 0.3375 ;
        RECT 1.8750 0.5625 1.9500 0.6375 ;
        RECT 1.4325 0.4350 1.5075 0.5100 ;
        RECT 1.3500 0.1650 1.4250 0.2400 ;
        RECT 1.1400 0.6600 1.2150 0.7350 ;
        RECT 0.9000 0.8025 0.9750 0.8775 ;
        RECT 0.2925 0.7125 0.3675 0.7875 ;
        LAYER M2 ;
        RECT 3.4125 0.2625 3.5175 0.6075 ;
        RECT 2.6625 0.2625 3.4125 0.3375 ;
        RECT 2.5875 0.2625 2.6625 0.8850 ;
        RECT 2.3700 0.7800 2.5875 0.8850 ;
        RECT 2.4300 0.3525 2.5050 0.5250 ;
        RECT 2.2950 0.6000 2.4675 0.6750 ;
        RECT 2.1450 0.4500 2.4300 0.5250 ;
        RECT 2.2200 0.6000 2.2950 0.9375 ;
        RECT 1.9950 0.2625 2.2800 0.3375 ;
        RECT 0.9750 0.8625 2.2200 0.9375 ;
        RECT 2.0700 0.4500 2.1450 0.7875 ;
        RECT 1.5075 0.7125 2.0700 0.7875 ;
        RECT 1.9200 0.2625 1.9950 0.6375 ;
        RECT 1.8150 0.5625 1.9200 0.6375 ;
        RECT 1.4325 0.3900 1.5075 0.7875 ;
        RECT 1.2600 0.1650 1.5000 0.2400 ;
        RECT 1.1850 0.1650 1.2600 0.7500 ;
        RECT 1.0950 0.6450 1.1850 0.7500 ;
        RECT 0.9000 0.7125 0.9750 0.9375 ;
        RECT 0.2475 0.7125 0.9000 0.7875 ;
    END
END DFCNQ_0111


MACRO DFCNQ_1010
    CLASS CORE ;
    FOREIGN DFCNQ_1010 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.9900 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 3.8775 0.2175 3.9525 0.8325 ;
        RECT 3.8475 0.2175 3.8775 0.3825 ;
        RECT 3.8475 0.6675 3.8775 0.8325 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.4500 0.5625 0.9150 0.6375 ;
        VIA 0.7125 0.6000 VIA12_square ;
        END
    END D
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.0675 0.4125 0.6225 0.4875 ;
        VIA 0.1800 0.4500 VIA12_square ;
        END
    END CP
    PIN CDN
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 3.4950 0.1125 3.5700 0.5775 ;
        RECT 1.7550 0.1125 3.4950 0.1875 ;
        RECT 1.6500 0.1125 1.7550 0.5250 ;
        VIA 3.5325 0.4875 VIA12_square ;
        VIA 1.7025 0.4425 VIA12_square ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 3.7350 -0.0750 3.9900 0.0750 ;
        RECT 3.6150 -0.0750 3.7350 0.1800 ;
        RECT 3.1050 -0.0750 3.6150 0.0750 ;
        RECT 2.9850 -0.0750 3.1050 0.2175 ;
        RECT 2.0550 -0.0750 2.9850 0.0750 ;
        RECT 1.9350 -0.0750 2.0550 0.1800 ;
        RECT 0.7875 -0.0750 1.9350 0.0750 ;
        RECT 0.6825 -0.0750 0.7875 0.2400 ;
        RECT 0.3750 -0.0750 0.6825 0.0750 ;
        RECT 0.2550 -0.0750 0.3750 0.1875 ;
        RECT 0.0000 -0.0750 0.2550 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 3.7350 0.9750 3.9900 1.1250 ;
        RECT 3.6150 0.8700 3.7350 1.1250 ;
        RECT 3.3000 0.9750 3.6150 1.1250 ;
        RECT 3.2250 0.8325 3.3000 1.1250 ;
        RECT 2.0550 0.9750 3.2250 1.1250 ;
        RECT 1.9500 0.8100 2.0550 1.1250 ;
        RECT 1.6350 0.9750 1.9500 1.1250 ;
        RECT 1.5150 0.8325 1.6350 1.1250 ;
        RECT 0.7725 0.9750 1.5150 1.1250 ;
        RECT 0.6975 0.7950 0.7725 1.1250 ;
        RECT 0.3750 0.9750 0.6975 1.1250 ;
        RECT 0.2550 0.8625 0.3750 1.1250 ;
        RECT 0.0000 0.9750 0.2550 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 3.8550 0.2700 3.9150 0.3300 ;
        RECT 3.8550 0.7200 3.9150 0.7800 ;
        RECT 3.7425 0.4950 3.8025 0.5550 ;
        RECT 3.6450 0.1200 3.7050 0.1800 ;
        RECT 3.6450 0.8700 3.7050 0.9300 ;
        RECT 3.5400 0.4725 3.6000 0.5325 ;
        RECT 3.4350 0.8325 3.4950 0.8925 ;
        RECT 3.3300 0.4950 3.3900 0.5550 ;
        RECT 3.2250 0.2775 3.2850 0.3375 ;
        RECT 3.2250 0.8625 3.2850 0.9225 ;
        RECT 3.1200 0.4950 3.1800 0.5550 ;
        RECT 3.0150 0.1575 3.0750 0.2175 ;
        RECT 3.0150 0.8325 3.0750 0.8925 ;
        RECT 2.9100 0.5100 2.9700 0.5700 ;
        RECT 2.7000 0.5250 2.7600 0.5850 ;
        RECT 2.5950 0.1725 2.6550 0.2325 ;
        RECT 2.5950 0.8325 2.6550 0.8925 ;
        RECT 2.4900 0.3750 2.5500 0.4350 ;
        RECT 2.3850 0.1725 2.4450 0.2325 ;
        RECT 2.3850 0.7350 2.4450 0.7950 ;
        RECT 2.2800 0.5175 2.3400 0.5775 ;
        RECT 2.1750 0.1575 2.2350 0.2175 ;
        RECT 2.1750 0.8175 2.2350 0.8775 ;
        RECT 2.0700 0.3750 2.1300 0.4350 ;
        RECT 1.9650 0.1200 2.0250 0.1800 ;
        RECT 1.9650 0.8400 2.0250 0.9000 ;
        RECT 1.8600 0.5400 1.9200 0.6000 ;
        RECT 1.7550 0.8325 1.8150 0.8925 ;
        RECT 1.6500 0.4800 1.7100 0.5400 ;
        RECT 1.5450 0.8325 1.6050 0.8925 ;
        RECT 1.4400 0.4575 1.5000 0.5175 ;
        RECT 1.3350 0.1800 1.3950 0.2400 ;
        RECT 1.3350 0.8100 1.3950 0.8700 ;
        RECT 1.2300 0.5025 1.2900 0.5625 ;
        RECT 1.1250 0.1725 1.1850 0.2325 ;
        RECT 1.1250 0.8025 1.1850 0.8625 ;
        RECT 1.0200 0.3600 1.0800 0.4200 ;
        RECT 0.9150 0.1725 0.9750 0.2325 ;
        RECT 0.8100 0.5250 0.8700 0.5850 ;
        RECT 0.7050 0.1575 0.7650 0.2175 ;
        RECT 0.7050 0.8325 0.7650 0.8925 ;
        RECT 0.4950 0.2775 0.5550 0.3375 ;
        RECT 0.4950 0.7350 0.5550 0.7950 ;
        RECT 0.3900 0.4650 0.4500 0.5250 ;
        RECT 0.2850 0.1200 0.3450 0.1800 ;
        RECT 0.2850 0.8700 0.3450 0.9300 ;
        RECT 0.1800 0.4875 0.2400 0.5475 ;
        RECT 0.0750 0.2400 0.1350 0.3000 ;
        RECT 0.0750 0.7500 0.1350 0.8100 ;
        LAYER M1 ;
        RECT 3.7575 0.4650 3.8025 0.5850 ;
        RECT 3.6825 0.2550 3.7575 0.7950 ;
        RECT 3.3900 0.2550 3.6825 0.3300 ;
        RECT 3.5400 0.7200 3.6825 0.7950 ;
        RECT 3.4725 0.4050 3.6075 0.6450 ;
        RECT 3.4650 0.7200 3.5400 0.9000 ;
        RECT 3.4050 0.8100 3.4650 0.9000 ;
        RECT 3.3225 0.2550 3.3900 0.3450 ;
        RECT 3.3150 0.4500 3.3900 0.7275 ;
        RECT 3.2400 0.2700 3.3225 0.3450 ;
        RECT 3.1425 0.6525 3.3150 0.7275 ;
        RECT 3.1650 0.2700 3.2400 0.5775 ;
        RECT 3.0150 0.4800 3.1650 0.5775 ;
        RECT 3.0825 0.6525 3.1425 0.7500 ;
        RECT 2.5500 0.8250 3.1200 0.9000 ;
        RECT 2.4450 0.6750 3.0825 0.7500 ;
        RECT 2.9100 0.4800 3.0150 0.6000 ;
        RECT 2.8800 0.3000 2.9700 0.4050 ;
        RECT 2.8050 0.1500 2.8800 0.4050 ;
        RECT 2.5725 0.1500 2.8050 0.2550 ;
        RECT 2.6775 0.5100 2.7900 0.5925 ;
        RECT 2.4150 0.3300 2.7150 0.4350 ;
        RECT 2.2500 0.5175 2.6775 0.5925 ;
        RECT 2.3400 0.1500 2.4675 0.2550 ;
        RECT 2.3700 0.6750 2.4450 0.8400 ;
        RECT 2.2350 0.1500 2.3400 0.4425 ;
        RECT 2.2125 0.8100 2.2650 0.8850 ;
        RECT 2.1450 0.1500 2.2350 0.2550 ;
        RECT 2.1375 0.6600 2.2125 0.8850 ;
        RECT 2.0475 0.3300 2.1600 0.4350 ;
        RECT 2.0250 0.6600 2.1375 0.7350 ;
        RECT 1.9725 0.2550 2.0475 0.4350 ;
        RECT 1.8600 0.5100 2.0250 0.7350 ;
        RECT 1.8450 0.2550 1.9725 0.3300 ;
        RECT 1.7700 0.1950 1.8450 0.3300 ;
        RECT 1.7850 0.8175 1.8450 0.9000 ;
        RECT 1.6200 0.4050 1.7850 0.6000 ;
        RECT 1.7100 0.6825 1.7850 0.9000 ;
        RECT 1.4850 0.1950 1.7700 0.2700 ;
        RECT 1.4400 0.6825 1.7100 0.7575 ;
        RECT 1.4250 0.3450 1.5300 0.6075 ;
        RECT 1.3350 0.1500 1.4850 0.2700 ;
        RECT 1.3350 0.6825 1.4400 0.9000 ;
        RECT 0.6000 0.3450 1.4250 0.4200 ;
        RECT 1.0200 0.4950 1.3200 0.5700 ;
        RECT 1.0950 0.6450 1.2600 0.9000 ;
        RECT 0.8925 0.1500 1.2300 0.2550 ;
        RECT 0.9450 0.4950 1.0200 0.9000 ;
        RECT 0.8550 0.7800 0.9450 0.9000 ;
        RECT 0.6750 0.4950 0.8700 0.6900 ;
        RECT 0.5625 0.2475 0.6000 0.7200 ;
        RECT 0.5250 0.2475 0.5625 0.8400 ;
        RECT 0.4875 0.2475 0.5250 0.3675 ;
        RECT 0.4875 0.6450 0.5250 0.8400 ;
        RECT 0.4125 0.4350 0.4500 0.5550 ;
        RECT 0.3375 0.2625 0.4125 0.7875 ;
        RECT 0.1425 0.2625 0.3375 0.3375 ;
        RECT 0.1425 0.7125 0.3375 0.7875 ;
        RECT 0.0975 0.4125 0.2625 0.6375 ;
        RECT 0.0675 0.2025 0.1425 0.3375 ;
        RECT 0.0675 0.7125 0.1425 0.8475 ;
        LAYER VIA1 ;
        RECT 2.8500 0.3225 2.9250 0.3975 ;
        RECT 2.8050 0.6750 2.8800 0.7500 ;
        RECT 2.6550 0.5175 2.7300 0.5925 ;
        RECT 2.4675 0.3450 2.5425 0.4200 ;
        RECT 2.2500 0.3300 2.3250 0.4050 ;
        RECT 1.9050 0.5100 1.9800 0.5850 ;
        RECT 1.4325 0.4875 1.5075 0.5625 ;
        RECT 1.3800 0.1950 1.4550 0.2700 ;
        RECT 1.1400 0.6600 1.2150 0.7350 ;
        RECT 0.9000 0.8025 0.9750 0.8775 ;
        RECT 0.2925 0.7125 0.3675 0.7875 ;
        LAYER M2 ;
        RECT 2.8800 0.3150 2.9700 0.4200 ;
        RECT 2.8050 0.3150 2.8800 0.7950 ;
        RECT 2.6550 0.4650 2.7300 0.8850 ;
        RECT 1.0200 0.8100 2.6550 0.8850 ;
        RECT 2.5125 0.3150 2.5800 0.4500 ;
        RECT 2.4375 0.3150 2.5125 0.7350 ;
        RECT 1.5075 0.6600 2.4375 0.7350 ;
        RECT 2.2125 0.3150 2.3625 0.4200 ;
        RECT 2.1375 0.3150 2.2125 0.5850 ;
        RECT 1.9650 0.5100 2.1375 0.5850 ;
        RECT 1.8600 0.4800 1.9650 0.5850 ;
        RECT 1.4325 0.4425 1.5075 0.7350 ;
        RECT 1.2600 0.1950 1.5000 0.2700 ;
        RECT 1.1850 0.1950 1.2600 0.7350 ;
        RECT 1.0950 0.6600 1.1850 0.7350 ;
        RECT 0.8550 0.7950 1.0200 0.8850 ;
        RECT 0.4650 0.7950 0.8550 0.8700 ;
        RECT 0.3900 0.7125 0.4650 0.8700 ;
        RECT 0.2475 0.7125 0.3900 0.7875 ;
    END
END DFCNQ_1010


MACRO DFCN_0011
    CLASS CORE ;
    FOREIGN DFCN_0011 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.6200 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 3.8175 0.2625 3.8925 0.7875 ;
        RECT 3.3600 0.2625 3.8175 0.3375 ;
        RECT 3.2775 0.7125 3.8175 0.7875 ;
        RECT 3.2550 0.2625 3.3600 0.4125 ;
        VIA 3.3900 0.7500 VIA12_square ;
        VIA 3.3075 0.3375 VIA12_square ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 4.5075 0.3075 4.5825 0.7425 ;
        RECT 4.3425 0.3075 4.5075 0.3825 ;
        RECT 4.3425 0.6675 4.5075 0.7425 ;
        RECT 4.2675 0.2175 4.3425 0.3825 ;
        RECT 4.2675 0.6675 4.3425 0.8325 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.4500 0.5625 0.9150 0.6375 ;
        VIA 0.7125 0.6000 VIA12_square ;
        END
    END D
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.0675 0.4125 0.6225 0.4875 ;
        VIA 0.1800 0.4500 VIA12_square ;
        END
    END CP
    PIN CDN
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 3.9675 0.1125 4.0425 0.6450 ;
        RECT 1.7550 0.1125 3.9675 0.1875 ;
        RECT 1.6800 0.1125 1.7550 0.4275 ;
        RECT 1.5825 0.3225 1.6800 0.4275 ;
        VIA 4.0050 0.5100 VIA12_square ;
        VIA 1.6725 0.3750 VIA12_square ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 4.5750 -0.0750 4.6200 0.0750 ;
        RECT 4.4550 -0.0750 4.5750 0.2325 ;
        RECT 4.1550 -0.0750 4.4550 0.0750 ;
        RECT 4.0350 -0.0750 4.1550 0.1800 ;
        RECT 3.5100 -0.0750 4.0350 0.0750 ;
        RECT 3.4350 -0.0750 3.5100 0.3000 ;
        RECT 3.0975 -0.0750 3.4350 0.0750 ;
        RECT 2.9925 -0.0750 3.0975 0.2925 ;
        RECT 2.0400 -0.0750 2.9925 0.0750 ;
        RECT 1.9650 -0.0750 2.0400 0.2550 ;
        RECT 0.7875 -0.0750 1.9650 0.0750 ;
        RECT 0.6825 -0.0750 0.7875 0.2400 ;
        RECT 0.3750 -0.0750 0.6825 0.0750 ;
        RECT 0.2550 -0.0750 0.3750 0.1875 ;
        RECT 0.0000 -0.0750 0.2550 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 4.5750 0.9750 4.6200 1.1250 ;
        RECT 4.4550 0.8175 4.5750 1.1250 ;
        RECT 4.1550 0.9750 4.4550 1.1250 ;
        RECT 4.0350 0.8625 4.1550 1.1250 ;
        RECT 3.5250 0.9750 4.0350 1.1250 ;
        RECT 3.4050 0.8625 3.5250 1.1250 ;
        RECT 3.1050 0.9750 3.4050 1.1250 ;
        RECT 2.9850 0.8700 3.1050 1.1250 ;
        RECT 2.0250 0.9750 2.9850 1.1250 ;
        RECT 1.9500 0.8400 2.0250 1.1250 ;
        RECT 1.6050 0.9750 1.9500 1.1250 ;
        RECT 1.5300 0.8025 1.6050 1.1250 ;
        RECT 0.7725 0.9750 1.5300 1.1250 ;
        RECT 0.6975 0.7950 0.7725 1.1250 ;
        RECT 0.3750 0.9750 0.6975 1.1250 ;
        RECT 0.2550 0.8625 0.3750 1.1250 ;
        RECT 0.0000 0.9750 0.2550 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 4.4850 0.1650 4.5450 0.2250 ;
        RECT 4.4850 0.8250 4.5450 0.8850 ;
        RECT 4.3725 0.4950 4.4325 0.5550 ;
        RECT 4.2750 0.2700 4.3350 0.3300 ;
        RECT 4.2750 0.7200 4.3350 0.7800 ;
        RECT 4.1700 0.4950 4.2300 0.5550 ;
        RECT 4.0650 0.1200 4.1250 0.1800 ;
        RECT 4.0650 0.8700 4.1250 0.9300 ;
        RECT 3.9600 0.4725 4.0200 0.5325 ;
        RECT 3.8550 0.7200 3.9150 0.7800 ;
        RECT 3.7425 0.4950 3.8025 0.5550 ;
        RECT 3.6450 0.1800 3.7050 0.2400 ;
        RECT 3.6450 0.7575 3.7050 0.8175 ;
        RECT 3.5400 0.4950 3.6000 0.5550 ;
        RECT 3.4350 0.2100 3.4950 0.2700 ;
        RECT 3.4350 0.8700 3.4950 0.9300 ;
        RECT 3.3225 0.4950 3.3825 0.5550 ;
        RECT 3.2250 0.2100 3.2850 0.2700 ;
        RECT 3.2250 0.7650 3.2850 0.8250 ;
        RECT 3.1200 0.4950 3.1800 0.5550 ;
        RECT 3.0150 0.2100 3.0750 0.2700 ;
        RECT 3.0150 0.8700 3.0750 0.9300 ;
        RECT 2.9025 0.5625 2.9625 0.6225 ;
        RECT 2.8050 0.1800 2.8650 0.2400 ;
        RECT 2.8050 0.8100 2.8650 0.8700 ;
        RECT 2.7000 0.5775 2.7600 0.6375 ;
        RECT 2.5950 0.1725 2.6550 0.2325 ;
        RECT 2.5950 0.8100 2.6550 0.8700 ;
        RECT 2.4900 0.4200 2.5500 0.4800 ;
        RECT 2.3850 0.1800 2.4450 0.2400 ;
        RECT 2.3850 0.8100 2.4450 0.8700 ;
        RECT 2.2875 0.5625 2.3475 0.6225 ;
        RECT 2.1750 0.1800 2.2350 0.2400 ;
        RECT 2.1750 0.8100 2.2350 0.8700 ;
        RECT 2.0625 0.4200 2.1225 0.4800 ;
        RECT 1.9650 0.1650 2.0250 0.2250 ;
        RECT 1.9650 0.8700 2.0250 0.9300 ;
        RECT 1.8600 0.5625 1.9200 0.6225 ;
        RECT 1.7550 0.8325 1.8150 0.8925 ;
        RECT 1.6500 0.4500 1.7100 0.5100 ;
        RECT 1.5450 0.8325 1.6050 0.8925 ;
        RECT 1.4400 0.4350 1.5000 0.4950 ;
        RECT 1.3350 0.1800 1.3950 0.2400 ;
        RECT 1.3350 0.8100 1.3950 0.8700 ;
        RECT 1.2225 0.5025 1.2825 0.5625 ;
        RECT 1.1250 0.1725 1.1850 0.2325 ;
        RECT 1.1250 0.8025 1.1850 0.8625 ;
        RECT 1.0200 0.3525 1.0800 0.4125 ;
        RECT 0.9150 0.1725 0.9750 0.2325 ;
        RECT 0.8100 0.5250 0.8700 0.5850 ;
        RECT 0.7050 0.1575 0.7650 0.2175 ;
        RECT 0.7050 0.8325 0.7650 0.8925 ;
        RECT 0.4950 0.2775 0.5550 0.3375 ;
        RECT 0.4950 0.7350 0.5550 0.7950 ;
        RECT 0.3900 0.4650 0.4500 0.5250 ;
        RECT 0.2850 0.1200 0.3450 0.1800 ;
        RECT 0.2850 0.8700 0.3450 0.9300 ;
        RECT 0.1800 0.4875 0.2400 0.5475 ;
        RECT 0.0750 0.2400 0.1350 0.3000 ;
        RECT 0.0750 0.7500 0.1350 0.8100 ;
        LAYER M1 ;
        RECT 4.1925 0.4650 4.4325 0.5850 ;
        RECT 4.1175 0.2625 4.1925 0.7875 ;
        RECT 3.9600 0.2625 4.1175 0.3375 ;
        RECT 3.7425 0.7125 4.1175 0.7875 ;
        RECT 3.8775 0.4125 4.0425 0.6150 ;
        RECT 3.8850 0.1500 3.9600 0.3375 ;
        RECT 3.6450 0.1500 3.8850 0.2700 ;
        RECT 3.5175 0.4575 3.8025 0.6075 ;
        RECT 3.6375 0.7125 3.7425 0.8475 ;
        RECT 3.3300 0.6825 3.5025 0.7875 ;
        RECT 3.1500 0.4875 3.4125 0.5625 ;
        RECT 3.2250 0.1500 3.3600 0.4125 ;
        RECT 3.2100 0.6825 3.3300 0.9000 ;
        RECT 3.0750 0.4125 3.1500 0.5625 ;
        RECT 3.0000 0.6375 3.1350 0.7950 ;
        RECT 2.9100 0.4125 3.0750 0.4875 ;
        RECT 2.9400 0.5625 3.0000 0.7950 ;
        RECT 2.8725 0.5625 2.9400 0.7050 ;
        RECT 2.8050 0.1500 2.9100 0.4875 ;
        RECT 2.5950 0.7800 2.8650 0.9000 ;
        RECT 2.2575 0.5625 2.7975 0.6750 ;
        RECT 2.6550 0.1500 2.7300 0.3825 ;
        RECT 2.5200 0.1500 2.6550 0.2850 ;
        RECT 2.3550 0.3600 2.5800 0.4875 ;
        RECT 2.3100 0.7500 2.5200 0.9000 ;
        RECT 2.2800 0.1500 2.4450 0.2700 ;
        RECT 2.2575 0.4125 2.3550 0.4875 ;
        RECT 2.1150 0.1500 2.2800 0.3375 ;
        RECT 2.1750 0.7800 2.2350 0.9000 ;
        RECT 2.1000 0.6600 2.1750 0.9000 ;
        RECT 1.8900 0.4125 2.1525 0.4875 ;
        RECT 1.9950 0.6600 2.1000 0.7350 ;
        RECT 1.8300 0.5625 1.9950 0.7350 ;
        RECT 1.8150 0.1500 1.8900 0.4875 ;
        RECT 1.7550 0.8175 1.8450 0.9000 ;
        RECT 1.4700 0.1500 1.8150 0.2250 ;
        RECT 1.6800 0.6225 1.7550 0.9000 ;
        RECT 1.5975 0.3000 1.7400 0.5475 ;
        RECT 1.4550 0.6225 1.6800 0.6975 ;
        RECT 1.4175 0.3450 1.5225 0.5475 ;
        RECT 1.3050 0.1500 1.4700 0.2700 ;
        RECT 1.3800 0.6225 1.4550 0.9000 ;
        RECT 0.6000 0.3450 1.4175 0.4200 ;
        RECT 1.3350 0.7575 1.3800 0.9000 ;
        RECT 1.0200 0.4950 1.3125 0.5700 ;
        RECT 1.0950 0.6450 1.2600 0.9000 ;
        RECT 0.8925 0.1500 1.2300 0.2550 ;
        RECT 0.9450 0.4950 1.0200 0.9000 ;
        RECT 0.8550 0.7800 0.9450 0.9000 ;
        RECT 0.6750 0.4950 0.8700 0.6900 ;
        RECT 0.5625 0.2475 0.6000 0.7200 ;
        RECT 0.5250 0.2475 0.5625 0.8400 ;
        RECT 0.4875 0.2475 0.5250 0.3675 ;
        RECT 0.4875 0.6450 0.5250 0.8400 ;
        RECT 0.4125 0.4350 0.4500 0.5550 ;
        RECT 0.3375 0.2625 0.4125 0.7875 ;
        RECT 0.1425 0.2625 0.3375 0.3375 ;
        RECT 0.1425 0.7125 0.3375 0.7875 ;
        RECT 0.0975 0.4125 0.2625 0.6375 ;
        RECT 0.0675 0.2025 0.1425 0.3375 ;
        RECT 0.0675 0.7125 0.1425 0.8475 ;
        LAYER VIA1 ;
        RECT 4.1175 0.6675 4.1925 0.7425 ;
        RECT 3.6375 0.5175 3.7125 0.5925 ;
        RECT 3.0075 0.7125 3.0825 0.7875 ;
        RECT 2.8800 0.4125 2.9550 0.4875 ;
        RECT 2.7375 0.8175 2.8125 0.8925 ;
        RECT 2.6550 0.2625 2.7300 0.3375 ;
        RECT 2.4300 0.3975 2.5050 0.4725 ;
        RECT 2.4075 0.7950 2.4825 0.8700 ;
        RECT 2.3175 0.6000 2.3925 0.6750 ;
        RECT 2.1600 0.2625 2.2350 0.3375 ;
        RECT 1.8750 0.5625 1.9500 0.6375 ;
        RECT 1.4325 0.4350 1.5075 0.5100 ;
        RECT 1.3500 0.1650 1.4250 0.2400 ;
        RECT 1.1400 0.6600 1.2150 0.7350 ;
        RECT 0.9000 0.8025 0.9750 0.8775 ;
        RECT 0.2925 0.7125 0.3675 0.7875 ;
        LAYER M2 ;
        RECT 4.1175 0.5550 4.1925 0.9375 ;
        RECT 3.1275 0.8625 4.1175 0.9375 ;
        RECT 3.6225 0.4800 3.7275 0.6375 ;
        RECT 3.1800 0.5625 3.6225 0.6375 ;
        RECT 3.1050 0.2625 3.1800 0.6375 ;
        RECT 3.0525 0.7125 3.1275 0.9375 ;
        RECT 2.6625 0.2625 3.1050 0.3375 ;
        RECT 2.9325 0.7125 3.0525 0.7875 ;
        RECT 2.9550 0.4125 3.0300 0.5325 ;
        RECT 2.8125 0.4125 2.9550 0.4875 ;
        RECT 2.8125 0.8625 2.9025 0.9375 ;
        RECT 2.7375 0.4125 2.8125 0.9375 ;
        RECT 2.5875 0.2625 2.6625 0.8850 ;
        RECT 2.3700 0.7800 2.5875 0.8850 ;
        RECT 2.4300 0.3525 2.5050 0.5250 ;
        RECT 2.2950 0.6000 2.4675 0.6750 ;
        RECT 2.1450 0.4500 2.4300 0.5250 ;
        RECT 2.2200 0.6000 2.2950 0.9375 ;
        RECT 1.9950 0.2625 2.2800 0.3375 ;
        RECT 0.9750 0.8625 2.2200 0.9375 ;
        RECT 2.0700 0.4500 2.1450 0.7875 ;
        RECT 1.5075 0.7125 2.0700 0.7875 ;
        RECT 1.9200 0.2625 1.9950 0.6375 ;
        RECT 1.8150 0.5625 1.9200 0.6375 ;
        RECT 1.4325 0.3900 1.5075 0.7875 ;
        RECT 1.2600 0.1650 1.5000 0.2400 ;
        RECT 1.1850 0.1650 1.2600 0.7500 ;
        RECT 1.0950 0.6450 1.1850 0.7500 ;
        RECT 0.9000 0.7125 0.9750 0.9375 ;
        RECT 0.2475 0.7125 0.9000 0.7875 ;
    END
END DFCN_0011


MACRO DFCN_0111
    CLASS CORE ;
    FOREIGN DFCN_0111 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.6700 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 4.9875 0.2400 5.3025 0.7650 ;
        VIA 5.1450 0.3225 VIA12_slot ;
        VIA 5.1450 0.6825 VIA12_slot ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 4.1475 0.2325 4.4625 0.7350 ;
        VIA 4.3050 0.3150 VIA12_slot ;
        VIA 4.3050 0.6525 VIA12_slot ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.4500 0.5625 0.9150 0.6375 ;
        VIA 0.7125 0.6000 VIA12_square ;
        END
    END D
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.0675 0.4125 0.6225 0.4875 ;
        VIA 0.1800 0.4500 VIA12_square ;
        END
    END CP
    PIN CDN
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 3.7275 0.1125 3.8025 0.7875 ;
        RECT 1.7550 0.1125 3.7275 0.1875 ;
        RECT 3.2550 0.7125 3.7275 0.7875 ;
        RECT 3.1800 0.4725 3.2550 0.7875 ;
        RECT 1.6800 0.1125 1.7550 0.4275 ;
        RECT 1.5825 0.3225 1.6800 0.4275 ;
        VIA 3.7650 0.5325 VIA12_square ;
        VIA 3.2175 0.5625 VIA12_square ;
        VIA 1.6725 0.3750 VIA12_square ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 5.6025 -0.0750 5.6700 0.0750 ;
        RECT 5.5275 -0.0750 5.6025 0.3225 ;
        RECT 5.2050 -0.0750 5.5275 0.0750 ;
        RECT 5.0850 -0.0750 5.2050 0.1950 ;
        RECT 4.7700 -0.0750 5.0850 0.0750 ;
        RECT 4.6950 -0.0750 4.7700 0.2850 ;
        RECT 4.3650 -0.0750 4.6950 0.0750 ;
        RECT 4.2450 -0.0750 4.3650 0.1875 ;
        RECT 3.9450 -0.0750 4.2450 0.0750 ;
        RECT 3.8400 -0.0750 3.9450 0.2250 ;
        RECT 3.0900 -0.0750 3.8400 0.0750 ;
        RECT 3.0000 -0.0750 3.0900 0.2625 ;
        RECT 2.0400 -0.0750 3.0000 0.0750 ;
        RECT 1.9650 -0.0750 2.0400 0.2550 ;
        RECT 0.7875 -0.0750 1.9650 0.0750 ;
        RECT 0.6825 -0.0750 0.7875 0.2400 ;
        RECT 0.3750 -0.0750 0.6825 0.0750 ;
        RECT 0.2550 -0.0750 0.3750 0.1875 ;
        RECT 0.0000 -0.0750 0.2550 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 5.6175 0.9750 5.6700 1.1250 ;
        RECT 5.5125 0.6450 5.6175 1.1250 ;
        RECT 5.2050 0.9750 5.5125 1.1250 ;
        RECT 5.0850 0.8175 5.2050 1.1250 ;
        RECT 4.7625 0.9750 5.0850 1.1250 ;
        RECT 4.6875 0.7500 4.7625 1.1250 ;
        RECT 4.3650 0.9750 4.6875 1.1250 ;
        RECT 4.2450 0.8175 4.3650 1.1250 ;
        RECT 3.9450 0.9750 4.2450 1.1250 ;
        RECT 3.8250 0.8700 3.9450 1.1250 ;
        RECT 3.5250 0.9750 3.8250 1.1250 ;
        RECT 3.4050 0.8700 3.5250 1.1250 ;
        RECT 3.1050 0.9750 3.4050 1.1250 ;
        RECT 2.9850 0.8700 3.1050 1.1250 ;
        RECT 2.0250 0.9750 2.9850 1.1250 ;
        RECT 1.9500 0.8400 2.0250 1.1250 ;
        RECT 1.6050 0.9750 1.9500 1.1250 ;
        RECT 1.5300 0.8025 1.6050 1.1250 ;
        RECT 0.7725 0.9750 1.5300 1.1250 ;
        RECT 0.6975 0.7950 0.7725 1.1250 ;
        RECT 0.3750 0.9750 0.6975 1.1250 ;
        RECT 0.2550 0.8625 0.3750 1.1250 ;
        RECT 0.0000 0.9750 0.2550 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 5.5350 0.2325 5.5950 0.2925 ;
        RECT 5.5350 0.6675 5.5950 0.7275 ;
        RECT 5.5350 0.8325 5.5950 0.8925 ;
        RECT 5.4300 0.4800 5.4900 0.5400 ;
        RECT 5.3250 0.2925 5.3850 0.3525 ;
        RECT 5.3250 0.6600 5.3850 0.7200 ;
        RECT 5.2200 0.4800 5.2800 0.5400 ;
        RECT 5.1150 0.1350 5.1750 0.1950 ;
        RECT 5.1150 0.8325 5.1750 0.8925 ;
        RECT 5.0100 0.4800 5.0700 0.5400 ;
        RECT 4.9050 0.2925 4.9650 0.3525 ;
        RECT 4.9050 0.6600 4.9650 0.7200 ;
        RECT 4.8000 0.4800 4.8600 0.5400 ;
        RECT 4.6950 0.1950 4.7550 0.2550 ;
        RECT 4.6950 0.7950 4.7550 0.8550 ;
        RECT 4.5900 0.4725 4.6500 0.5325 ;
        RECT 4.4850 0.2850 4.5450 0.3450 ;
        RECT 4.4850 0.6525 4.5450 0.7125 ;
        RECT 4.3800 0.4725 4.4400 0.5325 ;
        RECT 4.2750 0.1275 4.3350 0.1875 ;
        RECT 4.2750 0.8325 4.3350 0.8925 ;
        RECT 4.1700 0.4725 4.2300 0.5325 ;
        RECT 4.0650 0.2700 4.1250 0.3300 ;
        RECT 4.0650 0.6525 4.1250 0.7125 ;
        RECT 3.9600 0.4725 4.0200 0.5325 ;
        RECT 3.8550 0.1350 3.9150 0.1950 ;
        RECT 3.8550 0.8700 3.9150 0.9300 ;
        RECT 3.7500 0.4950 3.8100 0.5550 ;
        RECT 3.6450 0.1575 3.7050 0.2175 ;
        RECT 3.6450 0.7275 3.7050 0.7875 ;
        RECT 3.5400 0.4875 3.6000 0.5475 ;
        RECT 3.4350 0.3075 3.4950 0.3675 ;
        RECT 3.4350 0.8700 3.4950 0.9300 ;
        RECT 3.3375 0.4875 3.3975 0.5475 ;
        RECT 3.2250 0.1575 3.2850 0.2175 ;
        RECT 3.2250 0.7275 3.2850 0.7875 ;
        RECT 3.1200 0.4875 3.1800 0.5475 ;
        RECT 3.0150 0.1725 3.0750 0.2325 ;
        RECT 3.0150 0.8700 3.0750 0.9300 ;
        RECT 2.9100 0.5625 2.9700 0.6225 ;
        RECT 2.8050 0.1800 2.8650 0.2400 ;
        RECT 2.8050 0.8175 2.8650 0.8775 ;
        RECT 2.7000 0.5775 2.7600 0.6375 ;
        RECT 2.5950 0.1725 2.6550 0.2325 ;
        RECT 2.5950 0.8100 2.6550 0.8700 ;
        RECT 2.4900 0.4200 2.5500 0.4800 ;
        RECT 2.3850 0.1800 2.4450 0.2400 ;
        RECT 2.3850 0.8100 2.4450 0.8700 ;
        RECT 2.2875 0.5625 2.3475 0.6225 ;
        RECT 2.1750 0.1800 2.2350 0.2400 ;
        RECT 2.1750 0.8100 2.2350 0.8700 ;
        RECT 2.0625 0.4200 2.1225 0.4800 ;
        RECT 1.9650 0.1650 2.0250 0.2250 ;
        RECT 1.9650 0.8700 2.0250 0.9300 ;
        RECT 1.8600 0.5625 1.9200 0.6225 ;
        RECT 1.7550 0.8325 1.8150 0.8925 ;
        RECT 1.6500 0.4500 1.7100 0.5100 ;
        RECT 1.5450 0.8325 1.6050 0.8925 ;
        RECT 1.4400 0.4350 1.5000 0.4950 ;
        RECT 1.3350 0.1800 1.3950 0.2400 ;
        RECT 1.3350 0.8100 1.3950 0.8700 ;
        RECT 1.2225 0.5025 1.2825 0.5625 ;
        RECT 1.1250 0.1725 1.1850 0.2325 ;
        RECT 1.1250 0.8025 1.1850 0.8625 ;
        RECT 1.0200 0.3525 1.0800 0.4125 ;
        RECT 0.9150 0.1725 0.9750 0.2325 ;
        RECT 0.8100 0.5250 0.8700 0.5850 ;
        RECT 0.7050 0.1575 0.7650 0.2175 ;
        RECT 0.7050 0.8325 0.7650 0.8925 ;
        RECT 0.4950 0.2775 0.5550 0.3375 ;
        RECT 0.4950 0.7350 0.5550 0.7950 ;
        RECT 0.3900 0.4650 0.4500 0.5250 ;
        RECT 0.2850 0.1200 0.3450 0.1800 ;
        RECT 0.2850 0.8700 0.3450 0.9300 ;
        RECT 0.1800 0.4875 0.2400 0.5475 ;
        RECT 0.0750 0.2400 0.1350 0.3000 ;
        RECT 0.0750 0.7500 0.1350 0.8100 ;
        LAYER M1 ;
        RECT 4.7700 0.4575 5.5200 0.5625 ;
        RECT 4.8750 0.2700 5.4150 0.3675 ;
        RECT 4.8825 0.6375 5.4075 0.7425 ;
        RECT 4.5600 0.4350 4.6800 0.5400 ;
        RECT 4.1475 0.2625 4.5750 0.3600 ;
        RECT 4.0650 0.6150 4.5675 0.7425 ;
        RECT 3.9900 0.4650 4.5600 0.5400 ;
        RECT 4.0650 0.2400 4.1475 0.3600 ;
        RECT 3.9150 0.3000 3.9900 0.7950 ;
        RECT 3.3900 0.3000 3.9150 0.3750 ;
        RECT 3.0450 0.7200 3.9150 0.7950 ;
        RECT 3.6750 0.4500 3.8400 0.6450 ;
        RECT 3.1950 0.1500 3.7350 0.2250 ;
        RECT 3.3375 0.4500 3.6000 0.5775 ;
        RECT 3.1200 0.3675 3.2625 0.6450 ;
        RECT 2.9700 0.5625 3.0450 0.7950 ;
        RECT 2.9100 0.4125 3.0150 0.4875 ;
        RECT 2.8800 0.5625 2.9700 0.6675 ;
        RECT 2.8050 0.1500 2.9100 0.4875 ;
        RECT 2.5950 0.7800 2.8950 0.9000 ;
        RECT 2.2575 0.5625 2.7975 0.6750 ;
        RECT 2.6550 0.1500 2.7300 0.3825 ;
        RECT 2.5200 0.1500 2.6550 0.2850 ;
        RECT 2.3550 0.3600 2.5800 0.4875 ;
        RECT 2.3100 0.7500 2.5200 0.9000 ;
        RECT 2.2800 0.1500 2.4450 0.2700 ;
        RECT 2.2575 0.4125 2.3550 0.4875 ;
        RECT 2.1150 0.1500 2.2800 0.3375 ;
        RECT 2.1750 0.7800 2.2350 0.9000 ;
        RECT 2.1000 0.6600 2.1750 0.9000 ;
        RECT 1.8900 0.4125 2.1525 0.4875 ;
        RECT 1.9950 0.6600 2.1000 0.7350 ;
        RECT 1.8300 0.5625 1.9950 0.7350 ;
        RECT 1.8150 0.1500 1.8900 0.4875 ;
        RECT 1.7550 0.8175 1.8450 0.9000 ;
        RECT 1.4700 0.1500 1.8150 0.2250 ;
        RECT 1.6800 0.6225 1.7550 0.9000 ;
        RECT 1.5975 0.3000 1.7400 0.5475 ;
        RECT 1.4550 0.6225 1.6800 0.6975 ;
        RECT 1.4175 0.3450 1.5225 0.5475 ;
        RECT 1.3050 0.1500 1.4700 0.2700 ;
        RECT 1.3800 0.6225 1.4550 0.9000 ;
        RECT 0.6000 0.3450 1.4175 0.4200 ;
        RECT 1.3350 0.7575 1.3800 0.9000 ;
        RECT 1.0200 0.4950 1.3125 0.5700 ;
        RECT 1.0950 0.6450 1.2600 0.9000 ;
        RECT 0.8925 0.1500 1.2300 0.2550 ;
        RECT 0.9450 0.4950 1.0200 0.9000 ;
        RECT 0.8550 0.7800 0.9450 0.9000 ;
        RECT 0.6750 0.4950 0.8700 0.6900 ;
        RECT 0.5625 0.2475 0.6000 0.7200 ;
        RECT 0.5250 0.2475 0.5625 0.8400 ;
        RECT 0.4875 0.2475 0.5250 0.3675 ;
        RECT 0.4875 0.6450 0.5250 0.8400 ;
        RECT 0.4125 0.4350 0.4500 0.5550 ;
        RECT 0.3375 0.2625 0.4125 0.7875 ;
        RECT 0.1425 0.2625 0.3375 0.3375 ;
        RECT 0.1425 0.7125 0.3375 0.7875 ;
        RECT 0.0975 0.4125 0.2625 0.6375 ;
        RECT 0.0675 0.2025 0.1425 0.3375 ;
        RECT 0.0675 0.7125 0.1425 0.8475 ;
        LAYER VIA1 ;
        RECT 4.8150 0.4725 4.8900 0.5475 ;
        RECT 3.4275 0.4725 3.5025 0.5475 ;
        RECT 2.8500 0.4125 2.9250 0.4875 ;
        RECT 2.7375 0.8175 2.8125 0.8925 ;
        RECT 2.6550 0.2625 2.7300 0.3375 ;
        RECT 2.4300 0.3975 2.5050 0.4725 ;
        RECT 2.4075 0.7950 2.4825 0.8700 ;
        RECT 2.3175 0.6000 2.3925 0.6750 ;
        RECT 2.1600 0.2625 2.2350 0.3375 ;
        RECT 1.8750 0.5625 1.9500 0.6375 ;
        RECT 1.4325 0.4350 1.5075 0.5100 ;
        RECT 1.3500 0.1650 1.4250 0.2400 ;
        RECT 1.1400 0.6600 1.2150 0.7350 ;
        RECT 0.9000 0.8025 0.9750 0.8775 ;
        RECT 0.2925 0.7125 0.3675 0.7875 ;
        LAYER M2 ;
        RECT 4.7625 0.4275 4.9050 0.5925 ;
        RECT 4.6875 0.4275 4.7625 0.9375 ;
        RECT 2.8125 0.8625 4.6875 0.9375 ;
        RECT 3.4125 0.2625 3.5175 0.6075 ;
        RECT 2.6625 0.2625 3.4125 0.3375 ;
        RECT 2.8125 0.4125 3.0000 0.4875 ;
        RECT 2.7375 0.4125 2.8125 0.9375 ;
        RECT 2.5875 0.2625 2.6625 0.8850 ;
        RECT 2.3700 0.7800 2.5875 0.8850 ;
        RECT 2.4300 0.3525 2.5050 0.5250 ;
        RECT 2.2950 0.6000 2.4675 0.6750 ;
        RECT 2.1450 0.4500 2.4300 0.5250 ;
        RECT 2.2200 0.6000 2.2950 0.9375 ;
        RECT 1.9950 0.2625 2.2800 0.3375 ;
        RECT 0.9750 0.8625 2.2200 0.9375 ;
        RECT 2.0700 0.4500 2.1450 0.7875 ;
        RECT 1.5075 0.7125 2.0700 0.7875 ;
        RECT 1.9200 0.2625 1.9950 0.6375 ;
        RECT 1.8150 0.5625 1.9200 0.6375 ;
        RECT 1.4325 0.3900 1.5075 0.7875 ;
        RECT 1.2600 0.1650 1.5000 0.2400 ;
        RECT 1.1850 0.1650 1.2600 0.7500 ;
        RECT 1.0950 0.6450 1.1850 0.7500 ;
        RECT 0.9000 0.7125 0.9750 0.9375 ;
        RECT 0.2475 0.7125 0.9000 0.7875 ;
    END
END DFCN_0111


MACRO DFCN_1010
    CLASS CORE ;
    FOREIGN DFCN_1010 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.2000 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 3.1050 0.5625 3.5700 0.6375 ;
        VIA 3.2850 0.6000 VIA12_square ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 4.0875 0.2175 4.1625 0.8550 ;
        RECT 4.0575 0.2175 4.0875 0.3975 ;
        RECT 4.0575 0.6525 4.0875 0.8550 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.4500 0.5625 0.9150 0.6375 ;
        VIA 0.7125 0.6000 VIA12_square ;
        END
    END D
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.0675 0.4125 0.6225 0.4875 ;
        VIA 0.1800 0.4500 VIA12_square ;
        END
    END CP
    PIN CDN
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 3.7125 0.1125 3.7875 0.5775 ;
        RECT 1.7550 0.1125 3.7125 0.1875 ;
        RECT 1.6800 0.1125 1.7550 0.4275 ;
        RECT 1.5825 0.3225 1.6800 0.4275 ;
        VIA 3.7500 0.4650 VIA12_square ;
        VIA 1.6725 0.3750 VIA12_square ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 3.9450 -0.0750 4.2000 0.0750 ;
        RECT 3.8250 -0.0750 3.9450 0.1800 ;
        RECT 3.0975 -0.0750 3.8250 0.0750 ;
        RECT 2.9925 -0.0750 3.0975 0.2175 ;
        RECT 2.0400 -0.0750 2.9925 0.0750 ;
        RECT 1.9650 -0.0750 2.0400 0.2550 ;
        RECT 0.7875 -0.0750 1.9650 0.0750 ;
        RECT 0.6825 -0.0750 0.7875 0.2400 ;
        RECT 0.3750 -0.0750 0.6825 0.0750 ;
        RECT 0.2550 -0.0750 0.3750 0.1875 ;
        RECT 0.0000 -0.0750 0.2550 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 3.9450 0.9750 4.2000 1.1250 ;
        RECT 3.8250 0.8625 3.9450 1.1250 ;
        RECT 3.5100 0.9750 3.8250 1.1250 ;
        RECT 3.4050 0.8025 3.5100 1.1250 ;
        RECT 3.1050 0.9750 3.4050 1.1250 ;
        RECT 2.9850 0.8700 3.1050 1.1250 ;
        RECT 2.0250 0.9750 2.9850 1.1250 ;
        RECT 1.9500 0.8400 2.0250 1.1250 ;
        RECT 1.6050 0.9750 1.9500 1.1250 ;
        RECT 1.5300 0.8025 1.6050 1.1250 ;
        RECT 0.7725 0.9750 1.5300 1.1250 ;
        RECT 0.6975 0.7950 0.7725 1.1250 ;
        RECT 0.3750 0.9750 0.6975 1.1250 ;
        RECT 0.2550 0.8625 0.3750 1.1250 ;
        RECT 0.0000 0.9750 0.2550 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 4.0650 0.2625 4.1250 0.3225 ;
        RECT 4.0650 0.7425 4.1250 0.8025 ;
        RECT 3.9525 0.4950 4.0125 0.5550 ;
        RECT 3.8550 0.1200 3.9150 0.1800 ;
        RECT 3.8550 0.8700 3.9150 0.9300 ;
        RECT 3.7500 0.4725 3.8100 0.5325 ;
        RECT 3.6450 0.7875 3.7050 0.8475 ;
        RECT 3.5325 0.4950 3.5925 0.5550 ;
        RECT 3.4350 0.2475 3.4950 0.3075 ;
        RECT 3.4350 0.8325 3.4950 0.8925 ;
        RECT 3.2250 0.1725 3.2850 0.2325 ;
        RECT 3.2250 0.7350 3.2850 0.7950 ;
        RECT 3.1125 0.3975 3.1725 0.4575 ;
        RECT 3.0150 0.1350 3.0750 0.1950 ;
        RECT 3.0150 0.8700 3.0750 0.9300 ;
        RECT 2.9025 0.5625 2.9625 0.6225 ;
        RECT 2.8050 0.1800 2.8650 0.2400 ;
        RECT 2.8050 0.8175 2.8650 0.8775 ;
        RECT 2.7000 0.5775 2.7600 0.6375 ;
        RECT 2.5950 0.1725 2.6550 0.2325 ;
        RECT 2.5950 0.8100 2.6550 0.8700 ;
        RECT 2.4900 0.4200 2.5500 0.4800 ;
        RECT 2.3850 0.1800 2.4450 0.2400 ;
        RECT 2.3850 0.8100 2.4450 0.8700 ;
        RECT 2.2875 0.5625 2.3475 0.6225 ;
        RECT 2.1750 0.1800 2.2350 0.2400 ;
        RECT 2.1750 0.8100 2.2350 0.8700 ;
        RECT 2.0625 0.4200 2.1225 0.4800 ;
        RECT 1.9650 0.1650 2.0250 0.2250 ;
        RECT 1.9650 0.8700 2.0250 0.9300 ;
        RECT 1.8600 0.5625 1.9200 0.6225 ;
        RECT 1.7550 0.8325 1.8150 0.8925 ;
        RECT 1.6500 0.4500 1.7100 0.5100 ;
        RECT 1.5450 0.8325 1.6050 0.8925 ;
        RECT 1.4400 0.4350 1.5000 0.4950 ;
        RECT 1.3350 0.1800 1.3950 0.2400 ;
        RECT 1.3350 0.8100 1.3950 0.8700 ;
        RECT 1.2225 0.5025 1.2825 0.5625 ;
        RECT 1.1250 0.1725 1.1850 0.2325 ;
        RECT 1.1250 0.8025 1.1850 0.8625 ;
        RECT 1.0200 0.3525 1.0800 0.4125 ;
        RECT 0.9150 0.1725 0.9750 0.2325 ;
        RECT 0.8100 0.5250 0.8700 0.5850 ;
        RECT 0.7050 0.1575 0.7650 0.2175 ;
        RECT 0.7050 0.8325 0.7650 0.8925 ;
        RECT 0.4950 0.2775 0.5550 0.3375 ;
        RECT 0.4950 0.7350 0.5550 0.7950 ;
        RECT 0.3900 0.4650 0.4500 0.5250 ;
        RECT 0.2850 0.1200 0.3450 0.1800 ;
        RECT 0.2850 0.8700 0.3450 0.9300 ;
        RECT 0.1800 0.4875 0.2400 0.5475 ;
        RECT 0.0750 0.2400 0.1350 0.3000 ;
        RECT 0.0750 0.7500 0.1350 0.8100 ;
        LAYER M1 ;
        RECT 3.9825 0.4650 4.0125 0.5850 ;
        RECT 3.9075 0.2625 3.9825 0.7875 ;
        RECT 3.5100 0.2625 3.9075 0.3375 ;
        RECT 3.7350 0.7125 3.9075 0.7875 ;
        RECT 3.6675 0.4125 3.8325 0.6150 ;
        RECT 3.6150 0.7125 3.7350 0.8700 ;
        RECT 3.3975 0.4125 3.5925 0.6375 ;
        RECT 3.4200 0.2175 3.5100 0.3375 ;
        RECT 3.2475 0.1500 3.3225 0.8250 ;
        RECT 3.2025 0.1500 3.2475 0.2550 ;
        RECT 3.2175 0.7050 3.2475 0.8250 ;
        RECT 3.0825 0.3675 3.1725 0.4875 ;
        RECT 2.9700 0.5625 3.1425 0.7950 ;
        RECT 2.9100 0.4125 3.0825 0.4875 ;
        RECT 2.8725 0.5625 2.9700 0.6675 ;
        RECT 2.8050 0.1500 2.9100 0.4875 ;
        RECT 2.5950 0.7800 2.8950 0.9000 ;
        RECT 2.2575 0.5625 2.7975 0.6750 ;
        RECT 2.6550 0.1500 2.7300 0.3825 ;
        RECT 2.5200 0.1500 2.6550 0.2850 ;
        RECT 2.3550 0.3600 2.5800 0.4875 ;
        RECT 2.3100 0.7500 2.5200 0.9000 ;
        RECT 2.2800 0.1500 2.4450 0.2700 ;
        RECT 2.2575 0.4125 2.3550 0.4875 ;
        RECT 2.1150 0.1500 2.2800 0.3375 ;
        RECT 2.1750 0.7800 2.2350 0.9000 ;
        RECT 2.1000 0.6600 2.1750 0.9000 ;
        RECT 1.8900 0.4125 2.1525 0.4875 ;
        RECT 1.9950 0.6600 2.1000 0.7350 ;
        RECT 1.8300 0.5625 1.9950 0.7350 ;
        RECT 1.8150 0.1500 1.8900 0.4875 ;
        RECT 1.7550 0.8175 1.8450 0.9000 ;
        RECT 1.4700 0.1500 1.8150 0.2250 ;
        RECT 1.6800 0.6225 1.7550 0.9000 ;
        RECT 1.5975 0.3000 1.7400 0.5475 ;
        RECT 1.4550 0.6225 1.6800 0.6975 ;
        RECT 1.4175 0.3450 1.5225 0.5475 ;
        RECT 1.3050 0.1500 1.4700 0.2700 ;
        RECT 1.3800 0.6225 1.4550 0.9000 ;
        RECT 0.6000 0.3450 1.4175 0.4200 ;
        RECT 1.3350 0.7575 1.3800 0.9000 ;
        RECT 1.0200 0.4950 1.3125 0.5700 ;
        RECT 1.0950 0.6450 1.2600 0.9000 ;
        RECT 0.8925 0.1500 1.2300 0.2550 ;
        RECT 0.9450 0.4950 1.0200 0.9000 ;
        RECT 0.8550 0.7800 0.9450 0.9000 ;
        RECT 0.6750 0.4950 0.8700 0.6900 ;
        RECT 0.5625 0.2475 0.6000 0.7200 ;
        RECT 0.5250 0.2475 0.5625 0.8400 ;
        RECT 0.4875 0.2475 0.5250 0.3675 ;
        RECT 0.4875 0.6450 0.5250 0.8400 ;
        RECT 0.4125 0.4350 0.4500 0.5550 ;
        RECT 0.3375 0.2625 0.4125 0.7875 ;
        RECT 0.1425 0.2625 0.3375 0.3375 ;
        RECT 0.1425 0.7125 0.3375 0.7875 ;
        RECT 0.0975 0.4125 0.2625 0.6375 ;
        RECT 0.0675 0.2025 0.1425 0.3375 ;
        RECT 0.0675 0.7125 0.1425 0.8475 ;
        LAYER VIA1 ;
        RECT 3.6750 0.7125 3.7500 0.7875 ;
        RECT 3.4425 0.4125 3.5175 0.4875 ;
        RECT 3.0150 0.7125 3.0900 0.7875 ;
        RECT 2.8800 0.4125 2.9550 0.4875 ;
        RECT 2.7375 0.8175 2.8125 0.8925 ;
        RECT 2.6550 0.2625 2.7300 0.3375 ;
        RECT 2.4300 0.3975 2.5050 0.4725 ;
        RECT 2.4075 0.7950 2.4825 0.8700 ;
        RECT 2.3175 0.6000 2.3925 0.6750 ;
        RECT 2.1600 0.2625 2.2350 0.3375 ;
        RECT 1.8750 0.5625 1.9500 0.6375 ;
        RECT 1.4325 0.4350 1.5075 0.5100 ;
        RECT 1.3500 0.1650 1.4250 0.2400 ;
        RECT 1.1400 0.6600 1.2150 0.7350 ;
        RECT 0.9000 0.8025 0.9750 0.8775 ;
        RECT 0.2925 0.7125 0.3675 0.7875 ;
        LAYER M2 ;
        RECT 2.9400 0.7125 3.8250 0.7875 ;
        RECT 3.4275 0.4125 3.5625 0.4875 ;
        RECT 3.3525 0.2625 3.4275 0.4875 ;
        RECT 2.6625 0.2625 3.3525 0.3375 ;
        RECT 2.8125 0.4125 3.0300 0.4875 ;
        RECT 2.8125 0.8325 2.8425 0.9375 ;
        RECT 2.7375 0.4125 2.8125 0.9375 ;
        RECT 2.5875 0.2625 2.6625 0.8850 ;
        RECT 2.3700 0.7800 2.5875 0.8850 ;
        RECT 2.4300 0.3525 2.5050 0.5250 ;
        RECT 2.2950 0.6000 2.4675 0.6750 ;
        RECT 2.1450 0.4500 2.4300 0.5250 ;
        RECT 2.2200 0.6000 2.2950 0.9375 ;
        RECT 1.9950 0.2625 2.2800 0.3375 ;
        RECT 0.9750 0.8625 2.2200 0.9375 ;
        RECT 2.0700 0.4500 2.1450 0.7875 ;
        RECT 1.5075 0.7125 2.0700 0.7875 ;
        RECT 1.9200 0.2625 1.9950 0.6375 ;
        RECT 1.8150 0.5625 1.9200 0.6375 ;
        RECT 1.4325 0.3900 1.5075 0.7875 ;
        RECT 1.2600 0.1650 1.5000 0.2400 ;
        RECT 1.1850 0.1650 1.2600 0.7500 ;
        RECT 1.0950 0.6450 1.1850 0.7500 ;
        RECT 0.9000 0.7125 0.9750 0.9375 ;
        RECT 0.2475 0.7125 0.9000 0.7875 ;
    END
END DFCN_1010


MACRO DFQ_0011
    CLASS CORE ;
    FOREIGN DFQ_0011 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.5700 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 2.8050 0.2625 3.1950 0.3375 ;
        RECT 2.8050 0.7125 2.9400 0.7875 ;
        RECT 2.7300 0.2625 2.8050 0.7875 ;
        VIA 2.8575 0.3000 VIA12_square ;
        VIA 2.8575 0.7500 VIA12_square ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.3900 0.5625 0.8550 0.6375 ;
        VIA 0.7425 0.6000 VIA12_square ;
        END
    END D
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.0375 0.4125 0.2400 0.6375 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 3.3150 -0.0750 3.5700 0.0750 ;
        RECT 3.1950 -0.0750 3.3150 0.1875 ;
        RECT 2.8950 -0.0750 3.1950 0.0750 ;
        RECT 2.7750 -0.0750 2.8950 0.1875 ;
        RECT 1.8150 -0.0750 2.7750 0.0750 ;
        RECT 1.7100 -0.0750 1.8150 0.2100 ;
        RECT 0.7875 -0.0750 1.7100 0.0750 ;
        RECT 0.6825 -0.0750 0.7875 0.2400 ;
        RECT 0.3750 -0.0750 0.6825 0.0750 ;
        RECT 0.2550 -0.0750 0.3750 0.1875 ;
        RECT 0.0000 -0.0750 0.2550 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 3.3150 0.9750 3.5700 1.1250 ;
        RECT 3.1950 0.8625 3.3150 1.1250 ;
        RECT 2.8950 0.9750 3.1950 1.1250 ;
        RECT 2.7750 0.8625 2.8950 1.1250 ;
        RECT 1.8300 0.9750 2.7750 1.1250 ;
        RECT 1.7250 0.8250 1.8300 1.1250 ;
        RECT 0.7875 0.9750 1.7250 1.1250 ;
        RECT 0.6825 0.8100 0.7875 1.1250 ;
        RECT 0.3750 0.9750 0.6825 1.1250 ;
        RECT 0.2550 0.8625 0.3750 1.1250 ;
        RECT 0.0000 0.9750 0.2550 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 3.4350 0.2700 3.4950 0.3300 ;
        RECT 3.4350 0.8100 3.4950 0.8700 ;
        RECT 3.3225 0.4800 3.3825 0.5400 ;
        RECT 3.2250 0.1200 3.2850 0.1800 ;
        RECT 3.2250 0.8700 3.2850 0.9300 ;
        RECT 3.1200 0.4800 3.1800 0.5400 ;
        RECT 3.0150 0.2925 3.0750 0.3525 ;
        RECT 3.0150 0.6975 3.0750 0.7575 ;
        RECT 2.9100 0.4800 2.9700 0.5400 ;
        RECT 2.8050 0.1200 2.8650 0.1800 ;
        RECT 2.8050 0.8700 2.8650 0.9300 ;
        RECT 2.7000 0.4800 2.7600 0.5400 ;
        RECT 2.5950 0.8175 2.6550 0.8775 ;
        RECT 2.4900 0.3975 2.5500 0.4575 ;
        RECT 2.3850 0.1800 2.4450 0.2400 ;
        RECT 2.3850 0.8100 2.4450 0.8700 ;
        RECT 2.2800 0.5100 2.3400 0.5700 ;
        RECT 2.1750 0.1575 2.2350 0.2175 ;
        RECT 2.1750 0.8175 2.2350 0.8775 ;
        RECT 2.0700 0.3450 2.1300 0.4050 ;
        RECT 1.9650 0.1575 2.0250 0.2175 ;
        RECT 1.9650 0.8325 2.0250 0.8925 ;
        RECT 1.8525 0.6600 1.9125 0.7200 ;
        RECT 1.7550 0.1200 1.8150 0.1800 ;
        RECT 1.7550 0.8550 1.8150 0.9150 ;
        RECT 1.6575 0.3150 1.7175 0.3750 ;
        RECT 1.4400 0.3525 1.5000 0.4125 ;
        RECT 1.4400 0.6600 1.5000 0.7200 ;
        RECT 1.3350 0.1575 1.3950 0.2175 ;
        RECT 1.3350 0.8325 1.3950 0.8925 ;
        RECT 1.2300 0.3525 1.2900 0.4125 ;
        RECT 1.1250 0.1800 1.1850 0.2400 ;
        RECT 1.1250 0.8100 1.1850 0.8700 ;
        RECT 1.0200 0.5100 1.0800 0.5700 ;
        RECT 0.9150 0.8100 0.9750 0.8700 ;
        RECT 0.8100 0.5550 0.8700 0.6150 ;
        RECT 0.7050 0.1575 0.7650 0.2175 ;
        RECT 0.7050 0.8325 0.7650 0.8925 ;
        RECT 0.4950 0.2325 0.5550 0.2925 ;
        RECT 0.4950 0.7500 0.5550 0.8100 ;
        RECT 0.3900 0.4650 0.4500 0.5250 ;
        RECT 0.2850 0.1275 0.3450 0.1875 ;
        RECT 0.2850 0.8700 0.3450 0.9300 ;
        RECT 0.1800 0.4875 0.2400 0.5475 ;
        RECT 0.0750 0.2400 0.1350 0.3000 ;
        RECT 0.0750 0.7575 0.1350 0.8175 ;
        LAYER M1 ;
        RECT 3.4575 0.2625 3.5325 0.9000 ;
        RECT 3.2325 0.2625 3.4575 0.3375 ;
        RECT 3.4125 0.7800 3.4575 0.9000 ;
        RECT 3.3225 0.4425 3.3825 0.6975 ;
        RECT 3.3075 0.4425 3.3225 0.7875 ;
        RECT 3.1575 0.6225 3.3075 0.7875 ;
        RECT 3.1575 0.2625 3.2325 0.5475 ;
        RECT 2.6700 0.4725 3.1575 0.5475 ;
        RECT 2.7750 0.2625 3.0825 0.3825 ;
        RECT 2.7750 0.6675 3.0825 0.7875 ;
        RECT 2.3850 0.7725 2.7000 0.9000 ;
        RECT 2.3700 0.1500 2.6100 0.2850 ;
        RECT 2.4900 0.3600 2.5650 0.5025 ;
        RECT 2.2500 0.3600 2.4900 0.4350 ;
        RECT 2.1450 0.5100 2.4150 0.6300 ;
        RECT 2.1450 0.7050 2.3100 0.9000 ;
        RECT 1.9650 0.1500 2.2650 0.2250 ;
        RECT 2.1300 0.3000 2.2500 0.4350 ;
        RECT 2.0400 0.3000 2.1300 0.4050 ;
        RECT 1.9950 0.4800 2.0700 0.9000 ;
        RECT 1.9650 0.4800 1.9950 0.5550 ;
        RECT 1.9350 0.8250 1.9950 0.9000 ;
        RECT 1.8900 0.1500 1.9650 0.5550 ;
        RECT 1.8075 0.6300 1.9125 0.7500 ;
        RECT 1.6575 0.2850 1.8900 0.4050 ;
        RECT 1.6500 0.6675 1.8075 0.7500 ;
        RECT 1.5825 0.4800 1.7400 0.5925 ;
        RECT 1.5750 0.6675 1.6500 0.9000 ;
        RECT 1.5075 0.3450 1.5825 0.5550 ;
        RECT 1.3050 0.8250 1.5750 0.9000 ;
        RECT 0.6000 0.3450 1.5075 0.4200 ;
        RECT 1.4325 0.6300 1.5000 0.7500 ;
        RECT 1.0575 0.1500 1.4475 0.2550 ;
        RECT 1.3575 0.4950 1.4325 0.7500 ;
        RECT 0.9450 0.4950 1.3575 0.6000 ;
        RECT 0.8925 0.7800 1.1850 0.9000 ;
        RECT 0.6825 0.4950 0.8700 0.7050 ;
        RECT 0.5250 0.2025 0.6000 0.8325 ;
        RECT 0.4725 0.2025 0.5250 0.3225 ;
        RECT 0.4725 0.7275 0.5250 0.8325 ;
        RECT 0.3900 0.4275 0.4500 0.5625 ;
        RECT 0.3150 0.2625 0.3900 0.7875 ;
        RECT 0.1425 0.2625 0.3150 0.3375 ;
        RECT 0.1650 0.7125 0.3150 0.7875 ;
        RECT 0.0675 0.7125 0.1650 0.8700 ;
        RECT 0.0675 0.2025 0.1425 0.3375 ;
        LAYER VIA1 ;
        RECT 3.2025 0.7125 3.2775 0.7875 ;
        RECT 2.4300 0.1650 2.5050 0.2400 ;
        RECT 2.1900 0.5550 2.2650 0.6300 ;
        RECT 2.1900 0.8100 2.2650 0.8850 ;
        RECT 2.0925 0.3150 2.1675 0.3900 ;
        RECT 1.6275 0.5025 1.7025 0.5775 ;
        RECT 1.5750 0.7125 1.6500 0.7875 ;
        RECT 1.3200 0.5100 1.3950 0.5850 ;
        RECT 1.2000 0.1800 1.2750 0.2550 ;
        RECT 0.9900 0.5100 1.0650 0.5850 ;
        RECT 0.2700 0.7125 0.3450 0.7875 ;
        LAYER M2 ;
        RECT 3.1650 0.7125 3.3525 0.7875 ;
        RECT 3.0900 0.7125 3.1650 0.9375 ;
        RECT 2.5800 0.8625 3.0900 0.9375 ;
        RECT 2.5050 0.1650 2.5800 0.9375 ;
        RECT 2.3700 0.1650 2.5050 0.2400 ;
        RECT 2.1450 0.8100 2.5050 0.8850 ;
        RECT 1.7175 0.5550 2.3100 0.6300 ;
        RECT 2.0775 0.2625 2.1825 0.4350 ;
        RECT 1.5150 0.2625 2.0775 0.3375 ;
        RECT 1.6125 0.4650 1.7175 0.6300 ;
        RECT 1.2300 0.7125 1.6950 0.7875 ;
        RECT 1.4325 0.2625 1.5150 0.4200 ;
        RECT 1.4100 0.3450 1.4325 0.4200 ;
        RECT 1.3050 0.3450 1.4100 0.6225 ;
        RECT 1.2300 0.1650 1.3200 0.2700 ;
        RECT 1.1550 0.1650 1.2300 0.7875 ;
        RECT 0.9750 0.4650 1.0800 0.7875 ;
        RECT 0.2250 0.7125 0.9750 0.7875 ;
    END
END DFQ_0011


MACRO DFQ_0111
    CLASS CORE ;
    FOREIGN DFQ_0111 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.2000 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 3.5175 0.2400 3.8325 0.7650 ;
        VIA 3.6750 0.3225 VIA12_slot ;
        VIA 3.6750 0.6825 VIA12_slot ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.3900 0.5625 0.8550 0.6375 ;
        VIA 0.7425 0.6000 VIA12_square ;
        END
    END D
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.0375 0.4125 0.2400 0.6375 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 4.1325 -0.0750 4.2000 0.0750 ;
        RECT 4.0575 -0.0750 4.1325 0.3225 ;
        RECT 3.7350 -0.0750 4.0575 0.0750 ;
        RECT 3.6150 -0.0750 3.7350 0.1950 ;
        RECT 3.3075 -0.0750 3.6150 0.0750 ;
        RECT 3.2025 -0.0750 3.3075 0.2250 ;
        RECT 2.8950 -0.0750 3.2025 0.0750 ;
        RECT 2.7900 -0.0750 2.8950 0.2250 ;
        RECT 1.8150 -0.0750 2.7900 0.0750 ;
        RECT 1.7100 -0.0750 1.8150 0.2100 ;
        RECT 0.7875 -0.0750 1.7100 0.0750 ;
        RECT 0.6825 -0.0750 0.7875 0.2400 ;
        RECT 0.3750 -0.0750 0.6825 0.0750 ;
        RECT 0.2550 -0.0750 0.3750 0.1875 ;
        RECT 0.0000 -0.0750 0.2550 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 4.1475 0.9750 4.2000 1.1250 ;
        RECT 4.0425 0.6450 4.1475 1.1250 ;
        RECT 3.7350 0.9750 4.0425 1.1250 ;
        RECT 3.6150 0.8175 3.7350 1.1250 ;
        RECT 3.3075 0.9750 3.6150 1.1250 ;
        RECT 3.2025 0.8325 3.3075 1.1250 ;
        RECT 2.8725 0.9750 3.2025 1.1250 ;
        RECT 2.7975 0.8250 2.8725 1.1250 ;
        RECT 1.8300 0.9750 2.7975 1.1250 ;
        RECT 1.7250 0.8250 1.8300 1.1250 ;
        RECT 0.7875 0.9750 1.7250 1.1250 ;
        RECT 0.6825 0.8100 0.7875 1.1250 ;
        RECT 0.3750 0.9750 0.6825 1.1250 ;
        RECT 0.2550 0.8625 0.3750 1.1250 ;
        RECT 0.0000 0.9750 0.2550 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 4.0650 0.2325 4.1250 0.2925 ;
        RECT 4.0650 0.6675 4.1250 0.7275 ;
        RECT 4.0650 0.8325 4.1250 0.8925 ;
        RECT 3.9600 0.4800 4.0200 0.5400 ;
        RECT 3.8550 0.2925 3.9150 0.3525 ;
        RECT 3.8550 0.6600 3.9150 0.7200 ;
        RECT 3.7500 0.4800 3.8100 0.5400 ;
        RECT 3.6450 0.1350 3.7050 0.1950 ;
        RECT 3.6450 0.8325 3.7050 0.8925 ;
        RECT 3.5400 0.4800 3.6000 0.5400 ;
        RECT 3.4350 0.2925 3.4950 0.3525 ;
        RECT 3.4350 0.6600 3.4950 0.7200 ;
        RECT 3.3300 0.4800 3.3900 0.5400 ;
        RECT 3.2250 0.1425 3.2850 0.2025 ;
        RECT 3.2250 0.8550 3.2850 0.9150 ;
        RECT 3.1125 0.4875 3.1725 0.5475 ;
        RECT 3.0150 0.3000 3.0750 0.3600 ;
        RECT 3.0150 0.7200 3.0750 0.7800 ;
        RECT 2.9100 0.4950 2.9700 0.5550 ;
        RECT 2.8050 0.1350 2.8650 0.1950 ;
        RECT 2.8050 0.8550 2.8650 0.9150 ;
        RECT 2.7000 0.4575 2.7600 0.5175 ;
        RECT 2.5950 0.8175 2.6550 0.8775 ;
        RECT 2.4900 0.3975 2.5500 0.4575 ;
        RECT 2.3850 0.1800 2.4450 0.2400 ;
        RECT 2.3850 0.8100 2.4450 0.8700 ;
        RECT 2.2800 0.5100 2.3400 0.5700 ;
        RECT 2.1750 0.1575 2.2350 0.2175 ;
        RECT 2.1750 0.8175 2.2350 0.8775 ;
        RECT 2.0700 0.3450 2.1300 0.4050 ;
        RECT 1.9650 0.1575 2.0250 0.2175 ;
        RECT 1.9650 0.8325 2.0250 0.8925 ;
        RECT 1.8525 0.6600 1.9125 0.7200 ;
        RECT 1.7550 0.1200 1.8150 0.1800 ;
        RECT 1.7550 0.8550 1.8150 0.9150 ;
        RECT 1.6575 0.3150 1.7175 0.3750 ;
        RECT 1.4400 0.3525 1.5000 0.4125 ;
        RECT 1.4400 0.6600 1.5000 0.7200 ;
        RECT 1.3350 0.1575 1.3950 0.2175 ;
        RECT 1.3350 0.8325 1.3950 0.8925 ;
        RECT 1.2300 0.3525 1.2900 0.4125 ;
        RECT 1.1250 0.1800 1.1850 0.2400 ;
        RECT 1.1250 0.8100 1.1850 0.8700 ;
        RECT 1.0200 0.5100 1.0800 0.5700 ;
        RECT 0.9150 0.8100 0.9750 0.8700 ;
        RECT 0.8100 0.5250 0.8700 0.5850 ;
        RECT 0.7050 0.1575 0.7650 0.2175 ;
        RECT 0.7050 0.8325 0.7650 0.8925 ;
        RECT 0.4950 0.2325 0.5550 0.2925 ;
        RECT 0.4950 0.7500 0.5550 0.8100 ;
        RECT 0.3900 0.4650 0.4500 0.5250 ;
        RECT 0.2850 0.1275 0.3450 0.1875 ;
        RECT 0.2850 0.8700 0.3450 0.9300 ;
        RECT 0.1800 0.4875 0.2400 0.5475 ;
        RECT 0.0750 0.2400 0.1350 0.3000 ;
        RECT 0.0750 0.7575 0.1350 0.8175 ;
        LAYER M1 ;
        RECT 3.3300 0.4575 4.0500 0.5625 ;
        RECT 3.4050 0.2700 3.9450 0.3750 ;
        RECT 3.4125 0.6375 3.9375 0.7425 ;
        RECT 3.2550 0.3000 3.3300 0.7575 ;
        RECT 2.7600 0.3000 3.2550 0.3750 ;
        RECT 3.0825 0.6825 3.2550 0.7575 ;
        RECT 2.9100 0.4575 3.1725 0.5775 ;
        RECT 3.0075 0.6825 3.0825 0.8250 ;
        RECT 2.8350 0.4575 2.9100 0.6975 ;
        RECT 2.5200 0.6225 2.8350 0.6975 ;
        RECT 2.6850 0.3000 2.7600 0.5475 ;
        RECT 2.3850 0.7725 2.7000 0.9000 ;
        RECT 2.6550 0.4425 2.6850 0.5475 ;
        RECT 2.3700 0.1500 2.6100 0.2850 ;
        RECT 2.4900 0.3600 2.5650 0.5025 ;
        RECT 2.2500 0.3600 2.4900 0.4350 ;
        RECT 2.1450 0.5100 2.4150 0.6300 ;
        RECT 2.1450 0.7050 2.3100 0.9000 ;
        RECT 1.9650 0.1500 2.2650 0.2250 ;
        RECT 2.1300 0.3000 2.2500 0.4350 ;
        RECT 2.0400 0.3000 2.1300 0.4050 ;
        RECT 1.9950 0.4800 2.0700 0.9000 ;
        RECT 1.9650 0.4800 1.9950 0.5550 ;
        RECT 1.9350 0.8250 1.9950 0.9000 ;
        RECT 1.8900 0.1500 1.9650 0.5550 ;
        RECT 1.8075 0.6300 1.9125 0.7500 ;
        RECT 1.6575 0.2850 1.8900 0.4050 ;
        RECT 1.6500 0.6675 1.8075 0.7500 ;
        RECT 1.5825 0.4800 1.7400 0.5925 ;
        RECT 1.5750 0.6675 1.6500 0.9000 ;
        RECT 1.5075 0.3450 1.5825 0.5550 ;
        RECT 1.3050 0.8250 1.5750 0.9000 ;
        RECT 0.6000 0.3450 1.5075 0.4200 ;
        RECT 1.4325 0.6300 1.5000 0.7500 ;
        RECT 1.0575 0.1500 1.4475 0.2550 ;
        RECT 1.3575 0.4950 1.4325 0.7500 ;
        RECT 0.9450 0.4950 1.3575 0.6000 ;
        RECT 0.8925 0.7800 1.1850 0.9000 ;
        RECT 0.6825 0.4950 0.8700 0.7050 ;
        RECT 0.5250 0.2025 0.6000 0.8325 ;
        RECT 0.4725 0.2025 0.5250 0.3225 ;
        RECT 0.4725 0.7275 0.5250 0.8325 ;
        RECT 0.3900 0.4275 0.4500 0.5625 ;
        RECT 0.3150 0.2625 0.3900 0.7875 ;
        RECT 0.1425 0.2625 0.3150 0.3375 ;
        RECT 0.1650 0.7125 0.3150 0.7875 ;
        RECT 0.0675 0.7125 0.1650 0.8700 ;
        RECT 0.0675 0.2025 0.1425 0.3375 ;
        LAYER VIA1 ;
        RECT 2.5800 0.6225 2.6550 0.6975 ;
        RECT 2.4900 0.1650 2.5650 0.2400 ;
        RECT 2.1900 0.5550 2.2650 0.6300 ;
        RECT 2.1900 0.8100 2.2650 0.8850 ;
        RECT 2.0925 0.3150 2.1675 0.3900 ;
        RECT 1.6275 0.5025 1.7025 0.5775 ;
        RECT 1.5750 0.7125 1.6500 0.7875 ;
        RECT 1.3200 0.5100 1.3950 0.5850 ;
        RECT 1.2000 0.1800 1.2750 0.2550 ;
        RECT 0.9900 0.5100 1.0650 0.5850 ;
        RECT 0.2700 0.7125 0.3450 0.7875 ;
        LAYER M2 ;
        RECT 2.5800 0.1650 2.6550 0.8850 ;
        RECT 2.4300 0.1650 2.5800 0.2400 ;
        RECT 2.1450 0.8100 2.5800 0.8850 ;
        RECT 1.7175 0.5550 2.3100 0.6300 ;
        RECT 2.0775 0.2625 2.1825 0.4350 ;
        RECT 1.5150 0.2625 2.0775 0.3375 ;
        RECT 1.6125 0.4650 1.7175 0.6300 ;
        RECT 1.2300 0.7125 1.6950 0.7875 ;
        RECT 1.4325 0.2625 1.5150 0.4200 ;
        RECT 1.4100 0.3450 1.4325 0.4200 ;
        RECT 1.3050 0.3450 1.4100 0.6225 ;
        RECT 1.2300 0.1650 1.3200 0.2700 ;
        RECT 1.1550 0.1650 1.2300 0.7875 ;
        RECT 0.9750 0.4650 1.0800 0.7875 ;
        RECT 0.2250 0.7125 0.9750 0.7875 ;
    END
END DFQ_0111


MACRO DFQ_1010
    CLASS CORE ;
    FOREIGN DFQ_1010 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.5700 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 3.4575 0.2175 3.5325 0.8325 ;
        RECT 3.4275 0.2175 3.4575 0.3825 ;
        RECT 3.4275 0.6675 3.4575 0.8325 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.3900 0.5625 0.8550 0.6375 ;
        VIA 0.7425 0.6000 VIA12_square ;
        END
    END D
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.0375 0.4125 0.2400 0.6375 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 3.3075 -0.0750 3.5700 0.0750 ;
        RECT 3.2025 -0.0750 3.3075 0.3000 ;
        RECT 2.8875 -0.0750 3.2025 0.0750 ;
        RECT 2.7825 -0.0750 2.8875 0.2250 ;
        RECT 1.8150 -0.0750 2.7825 0.0750 ;
        RECT 1.7100 -0.0750 1.8150 0.2100 ;
        RECT 0.7875 -0.0750 1.7100 0.0750 ;
        RECT 0.6825 -0.0750 0.7875 0.2400 ;
        RECT 0.3750 -0.0750 0.6825 0.0750 ;
        RECT 0.2550 -0.0750 0.3750 0.1875 ;
        RECT 0.0000 -0.0750 0.2550 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 3.3075 0.9750 3.5700 1.1250 ;
        RECT 3.2025 0.6450 3.3075 1.1250 ;
        RECT 2.8875 0.9750 3.2025 1.1250 ;
        RECT 2.7825 0.8175 2.8875 1.1250 ;
        RECT 1.8300 0.9750 2.7825 1.1250 ;
        RECT 1.7250 0.8250 1.8300 1.1250 ;
        RECT 0.7875 0.9750 1.7250 1.1250 ;
        RECT 0.6825 0.8100 0.7875 1.1250 ;
        RECT 0.3750 0.9750 0.6825 1.1250 ;
        RECT 0.2550 0.8625 0.3750 1.1250 ;
        RECT 0.0000 0.9750 0.2550 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 3.4350 0.2700 3.4950 0.3300 ;
        RECT 3.4350 0.7200 3.4950 0.7800 ;
        RECT 3.3225 0.4725 3.3825 0.5325 ;
        RECT 3.2250 0.2175 3.2850 0.2775 ;
        RECT 3.2250 0.6675 3.2850 0.7275 ;
        RECT 3.2250 0.8325 3.2850 0.8925 ;
        RECT 3.0150 0.3000 3.0750 0.3600 ;
        RECT 3.0150 0.8100 3.0750 0.8700 ;
        RECT 2.9100 0.4875 2.9700 0.5475 ;
        RECT 2.8050 0.1425 2.8650 0.2025 ;
        RECT 2.8050 0.8550 2.8650 0.9150 ;
        RECT 2.7000 0.4725 2.7600 0.5325 ;
        RECT 2.5950 0.8175 2.6550 0.8775 ;
        RECT 2.4900 0.4950 2.5500 0.5550 ;
        RECT 2.3850 0.1800 2.4450 0.2400 ;
        RECT 2.3850 0.8100 2.4450 0.8700 ;
        RECT 2.2800 0.5100 2.3400 0.5700 ;
        RECT 2.1750 0.1575 2.2350 0.2175 ;
        RECT 2.1750 0.8175 2.2350 0.8775 ;
        RECT 2.0700 0.3450 2.1300 0.4050 ;
        RECT 1.9650 0.1575 2.0250 0.2175 ;
        RECT 1.9650 0.8325 2.0250 0.8925 ;
        RECT 1.8600 0.6600 1.9200 0.7200 ;
        RECT 1.7550 0.1200 1.8150 0.1800 ;
        RECT 1.7550 0.8550 1.8150 0.9150 ;
        RECT 1.6575 0.3150 1.7175 0.3750 ;
        RECT 1.4400 0.3525 1.5000 0.4125 ;
        RECT 1.4400 0.6600 1.5000 0.7200 ;
        RECT 1.3350 0.1575 1.3950 0.2175 ;
        RECT 1.3350 0.8325 1.3950 0.8925 ;
        RECT 1.2300 0.3525 1.2900 0.4125 ;
        RECT 1.1250 0.1800 1.1850 0.2400 ;
        RECT 1.1250 0.8100 1.1850 0.8700 ;
        RECT 1.0200 0.5100 1.0800 0.5700 ;
        RECT 0.9150 0.8100 0.9750 0.8700 ;
        RECT 0.8100 0.5250 0.8700 0.5850 ;
        RECT 0.7050 0.1575 0.7650 0.2175 ;
        RECT 0.7050 0.8325 0.7650 0.8925 ;
        RECT 0.4950 0.2325 0.5550 0.2925 ;
        RECT 0.4950 0.7500 0.5550 0.8100 ;
        RECT 0.3900 0.4650 0.4500 0.5250 ;
        RECT 0.2850 0.1275 0.3450 0.1875 ;
        RECT 0.2850 0.8700 0.3450 0.9300 ;
        RECT 0.1800 0.4875 0.2400 0.5475 ;
        RECT 0.0750 0.2400 0.1350 0.3000 ;
        RECT 0.0750 0.7575 0.1350 0.8175 ;
        LAYER M1 ;
        RECT 3.1275 0.4425 3.3825 0.5625 ;
        RECT 3.0525 0.3000 3.1275 0.9000 ;
        RECT 2.7600 0.3000 3.0525 0.3750 ;
        RECT 2.9925 0.7800 3.0525 0.9000 ;
        RECT 2.8350 0.4500 2.9775 0.7050 ;
        RECT 2.6850 0.3000 2.7600 0.5700 ;
        RECT 2.3850 0.7725 2.7000 0.9000 ;
        RECT 2.3700 0.1500 2.6100 0.2850 ;
        RECT 2.4900 0.3600 2.6100 0.5925 ;
        RECT 2.2500 0.3600 2.4900 0.4350 ;
        RECT 2.1450 0.5100 2.4150 0.6300 ;
        RECT 2.1450 0.7050 2.3100 0.9000 ;
        RECT 1.9650 0.1500 2.2650 0.2250 ;
        RECT 2.1300 0.3000 2.2500 0.4350 ;
        RECT 2.0400 0.3000 2.1300 0.4050 ;
        RECT 1.9950 0.4800 2.0700 0.9000 ;
        RECT 1.9650 0.4800 1.9950 0.5550 ;
        RECT 1.9350 0.8250 1.9950 0.9000 ;
        RECT 1.8900 0.1500 1.9650 0.5550 ;
        RECT 1.8075 0.6300 1.9200 0.7500 ;
        RECT 1.6575 0.2850 1.8900 0.4050 ;
        RECT 1.6500 0.6675 1.8075 0.7500 ;
        RECT 1.5825 0.4800 1.7400 0.5925 ;
        RECT 1.5750 0.6675 1.6500 0.9000 ;
        RECT 1.5075 0.3450 1.5825 0.5550 ;
        RECT 1.3050 0.8250 1.5750 0.9000 ;
        RECT 0.6000 0.3450 1.5075 0.4200 ;
        RECT 1.4325 0.6300 1.5000 0.7500 ;
        RECT 1.0575 0.1500 1.4475 0.2550 ;
        RECT 1.3575 0.4950 1.4325 0.7500 ;
        RECT 0.9450 0.4950 1.3575 0.6000 ;
        RECT 0.8925 0.7800 1.1850 0.9000 ;
        RECT 0.6825 0.4950 0.8700 0.7050 ;
        RECT 0.5250 0.2025 0.6000 0.8325 ;
        RECT 0.4725 0.2025 0.5250 0.3225 ;
        RECT 0.4725 0.7275 0.5250 0.8325 ;
        RECT 0.3900 0.4275 0.4500 0.5625 ;
        RECT 0.3150 0.2625 0.3900 0.7875 ;
        RECT 0.1425 0.2625 0.3150 0.3375 ;
        RECT 0.1650 0.7125 0.3150 0.7875 ;
        RECT 0.0675 0.7125 0.1650 0.8700 ;
        RECT 0.0675 0.2025 0.1425 0.3375 ;
        LAYER VIA1 ;
        RECT 2.8500 0.5625 2.9250 0.6375 ;
        RECT 2.4075 0.1650 2.4825 0.2400 ;
        RECT 2.1900 0.5175 2.2650 0.5925 ;
        RECT 2.1900 0.7125 2.2650 0.7875 ;
        RECT 2.0925 0.3150 2.1675 0.3900 ;
        RECT 1.6275 0.5025 1.7025 0.5775 ;
        RECT 1.5750 0.7125 1.6500 0.7875 ;
        RECT 1.3200 0.5100 1.3950 0.5850 ;
        RECT 1.2000 0.1800 1.2750 0.2550 ;
        RECT 0.9900 0.5100 1.0650 0.5850 ;
        RECT 0.2700 0.7125 0.3450 0.7875 ;
        LAYER M2 ;
        RECT 2.5350 0.5625 3.0000 0.6375 ;
        RECT 2.4600 0.1650 2.5350 0.7875 ;
        RECT 2.3475 0.1650 2.4600 0.2400 ;
        RECT 2.1450 0.7125 2.4600 0.7875 ;
        RECT 1.7475 0.5175 2.3100 0.5925 ;
        RECT 2.0775 0.2625 2.1825 0.4350 ;
        RECT 1.5150 0.2625 2.0775 0.3375 ;
        RECT 1.5825 0.4875 1.7475 0.5925 ;
        RECT 1.2300 0.7125 1.6950 0.7875 ;
        RECT 1.4325 0.2625 1.5150 0.4200 ;
        RECT 1.4100 0.3450 1.4325 0.4200 ;
        RECT 1.3050 0.3450 1.4100 0.6225 ;
        RECT 1.2300 0.1650 1.3200 0.2700 ;
        RECT 1.1550 0.1650 1.2300 0.7875 ;
        RECT 0.9750 0.4650 1.0800 0.7875 ;
        RECT 0.2250 0.7125 0.9750 0.7875 ;
    END
END DFQ_1010


MACRO DFSNQ_0011
    CLASS CORE ;
    FOREIGN DFSNQ_0011 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.2000 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN SDN
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 3.1575 0.4125 3.3000 0.4875 ;
        RECT 3.0825 0.4125 3.1575 0.9375 ;
        RECT 2.4525 0.8625 3.0825 0.9375 ;
        RECT 2.3775 0.5025 2.4525 0.9375 ;
        RECT 2.2350 0.5025 2.3775 0.6075 ;
        VIA 3.1875 0.4500 VIA12_square ;
        VIA 2.3175 0.5550 VIA12_square ;
        END
    END SDN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 3.6075 0.2625 3.6825 0.7125 ;
        RECT 3.1275 0.2625 3.6075 0.3375 ;
        RECT 3.4875 0.6375 3.6075 0.7125 ;
        VIA 3.6450 0.3600 VIA12_square ;
        VIA 3.6000 0.6750 VIA12_square ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.3900 0.5625 0.8550 0.6375 ;
        VIA 0.7425 0.6000 VIA12_square ;
        END
    END D
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.0375 0.4125 0.2400 0.6375 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 3.9450 -0.0750 4.2000 0.0750 ;
        RECT 3.8250 -0.0750 3.9450 0.2175 ;
        RECT 3.5175 -0.0750 3.8250 0.0750 ;
        RECT 3.4125 -0.0750 3.5175 0.2175 ;
        RECT 2.0550 -0.0750 3.4125 0.0750 ;
        RECT 1.9350 -0.0750 2.0550 0.2250 ;
        RECT 1.8450 -0.0750 1.9350 0.0750 ;
        RECT 1.7250 -0.0750 1.8450 0.2250 ;
        RECT 0.7875 -0.0750 1.7250 0.0750 ;
        RECT 0.6825 -0.0750 0.7875 0.2400 ;
        RECT 0.3750 -0.0750 0.6825 0.0750 ;
        RECT 0.2550 -0.0750 0.3750 0.1875 ;
        RECT 0.0000 -0.0750 0.2550 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 3.9450 0.9750 4.2000 1.1250 ;
        RECT 3.8250 0.8625 3.9450 1.1250 ;
        RECT 3.5175 0.9750 3.8250 1.1250 ;
        RECT 3.4125 0.8025 3.5175 1.1250 ;
        RECT 3.1050 0.9750 3.4125 1.1250 ;
        RECT 2.9850 0.8325 3.1050 1.1250 ;
        RECT 2.2650 0.9750 2.9850 1.1250 ;
        RECT 2.1450 0.8325 2.2650 1.1250 ;
        RECT 1.8450 0.9750 2.1450 1.1250 ;
        RECT 1.7250 0.8400 1.8450 1.1250 ;
        RECT 0.7875 0.9750 1.7250 1.1250 ;
        RECT 0.6825 0.8100 0.7875 1.1250 ;
        RECT 0.3750 0.9750 0.6825 1.1250 ;
        RECT 0.2550 0.8625 0.3750 1.1250 ;
        RECT 0.0000 0.9750 0.2550 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 4.0650 0.1800 4.1250 0.2400 ;
        RECT 4.0650 0.7200 4.1250 0.7800 ;
        RECT 3.9525 0.4950 4.0125 0.5550 ;
        RECT 3.8550 0.1425 3.9150 0.2025 ;
        RECT 3.8550 0.8625 3.9150 0.9225 ;
        RECT 3.7500 0.4950 3.8100 0.5550 ;
        RECT 3.6450 0.2325 3.7050 0.2925 ;
        RECT 3.6450 0.7350 3.7050 0.7950 ;
        RECT 3.5400 0.4950 3.6000 0.5550 ;
        RECT 3.4350 0.1275 3.4950 0.1875 ;
        RECT 3.4350 0.8325 3.4950 0.8925 ;
        RECT 3.3300 0.4725 3.3900 0.5325 ;
        RECT 3.2250 0.8025 3.2850 0.8625 ;
        RECT 3.1200 0.4800 3.1800 0.5400 ;
        RECT 3.0150 0.8325 3.0750 0.8925 ;
        RECT 2.9100 0.5175 2.9700 0.5775 ;
        RECT 2.8050 0.1800 2.8650 0.2400 ;
        RECT 2.8050 0.8100 2.8650 0.8700 ;
        RECT 2.7000 0.3600 2.7600 0.4200 ;
        RECT 2.5950 0.1725 2.6550 0.2325 ;
        RECT 2.5950 0.7650 2.6550 0.8250 ;
        RECT 2.4900 0.4950 2.5500 0.5550 ;
        RECT 2.3850 0.1725 2.4450 0.2325 ;
        RECT 2.3850 0.8025 2.4450 0.8625 ;
        RECT 2.2800 0.5100 2.3400 0.5700 ;
        RECT 2.1750 0.8325 2.2350 0.8925 ;
        RECT 2.0625 0.5100 2.1225 0.5700 ;
        RECT 1.9650 0.1575 2.0250 0.2175 ;
        RECT 1.9650 0.6900 2.0250 0.7500 ;
        RECT 1.8600 0.5100 1.9200 0.5700 ;
        RECT 1.7550 0.1575 1.8150 0.2175 ;
        RECT 1.7550 0.8475 1.8150 0.9075 ;
        RECT 1.6500 0.5100 1.7100 0.5700 ;
        RECT 1.4400 0.3450 1.5000 0.4050 ;
        RECT 1.4400 0.6450 1.5000 0.7050 ;
        RECT 1.3350 0.1575 1.3950 0.2175 ;
        RECT 1.3350 0.8250 1.3950 0.8850 ;
        RECT 1.2300 0.3450 1.2900 0.4050 ;
        RECT 1.1250 0.1575 1.1850 0.2175 ;
        RECT 1.1250 0.8100 1.1850 0.8700 ;
        RECT 1.0200 0.5025 1.0800 0.5625 ;
        RECT 0.9150 0.8100 0.9750 0.8700 ;
        RECT 0.8100 0.4950 0.8700 0.5550 ;
        RECT 0.7050 0.1575 0.7650 0.2175 ;
        RECT 0.7050 0.8325 0.7650 0.8925 ;
        RECT 0.4950 0.2325 0.5550 0.2925 ;
        RECT 0.4950 0.7500 0.5550 0.8100 ;
        RECT 0.3900 0.4650 0.4500 0.5250 ;
        RECT 0.2850 0.1275 0.3450 0.1875 ;
        RECT 0.2850 0.8700 0.3450 0.9300 ;
        RECT 0.1800 0.4875 0.2400 0.5475 ;
        RECT 0.0750 0.2400 0.1350 0.3000 ;
        RECT 0.0750 0.7575 0.1350 0.8175 ;
        LAYER M1 ;
        RECT 4.0875 0.1500 4.1625 0.7875 ;
        RECT 4.0575 0.1500 4.0875 0.2700 ;
        RECT 3.8625 0.7125 4.0875 0.7875 ;
        RECT 3.9375 0.3300 4.0125 0.5925 ;
        RECT 3.8025 0.2925 3.9375 0.4125 ;
        RECT 3.7875 0.4875 3.8625 0.7875 ;
        RECT 3.4350 0.4875 3.7875 0.5625 ;
        RECT 3.6000 0.1500 3.7275 0.4125 ;
        RECT 3.6075 0.6375 3.7125 0.8700 ;
        RECT 3.4875 0.6375 3.6075 0.7125 ;
        RECT 3.5100 0.3075 3.6000 0.4125 ;
        RECT 3.3300 0.4425 3.4350 0.5625 ;
        RECT 3.2025 0.6825 3.3150 0.8925 ;
        RECT 2.9175 0.1500 3.2625 0.2550 ;
        RECT 3.1050 0.3450 3.2550 0.6075 ;
        RECT 2.9100 0.6825 3.2025 0.7575 ;
        RECT 2.5950 0.4950 3.0000 0.5850 ;
        RECT 2.8050 0.1500 2.9175 0.2700 ;
        RECT 2.8050 0.6825 2.9100 0.9000 ;
        RECT 2.7375 0.3450 2.8200 0.4200 ;
        RECT 2.6700 0.3075 2.7375 0.4200 ;
        RECT 2.5200 0.6600 2.7300 0.8700 ;
        RECT 2.2050 0.1500 2.6850 0.2325 ;
        RECT 1.8000 0.3075 2.6700 0.3825 ;
        RECT 2.4900 0.4650 2.5950 0.5850 ;
        RECT 2.3400 0.6825 2.4450 0.8925 ;
        RECT 2.2050 0.4575 2.4150 0.6075 ;
        RECT 1.7250 0.6825 2.3400 0.7575 ;
        RECT 1.8000 0.4800 2.1225 0.6000 ;
        RECT 1.7250 0.3075 1.8000 0.4050 ;
        RECT 0.6000 0.3300 1.7250 0.4050 ;
        RECT 1.6500 0.4800 1.7250 0.7575 ;
        RECT 1.5750 0.4800 1.6500 0.6375 ;
        RECT 1.2900 0.8100 1.5900 0.9000 ;
        RECT 1.4175 0.6150 1.5000 0.7350 ;
        RECT 1.0800 0.1500 1.4400 0.2550 ;
        RECT 1.3425 0.4950 1.4175 0.7350 ;
        RECT 0.9825 0.4950 1.3425 0.6000 ;
        RECT 0.8925 0.7800 1.1850 0.9000 ;
        RECT 0.6825 0.4800 0.9075 0.7050 ;
        RECT 0.5250 0.2025 0.6000 0.8325 ;
        RECT 0.4725 0.2025 0.5250 0.3225 ;
        RECT 0.4725 0.7275 0.5250 0.8325 ;
        RECT 0.3900 0.4275 0.4500 0.5625 ;
        RECT 0.3150 0.2625 0.3900 0.7875 ;
        RECT 0.1425 0.2625 0.3150 0.3375 ;
        RECT 0.1650 0.7125 0.3150 0.7875 ;
        RECT 0.0675 0.7125 0.1650 0.8700 ;
        RECT 0.0675 0.2025 0.1425 0.3375 ;
        LAYER VIA1 ;
        RECT 3.9375 0.4125 4.0125 0.4875 ;
        RECT 2.9325 0.1650 3.0075 0.2400 ;
        RECT 2.7450 0.4950 2.8200 0.5700 ;
        RECT 2.5875 0.6600 2.6625 0.7350 ;
        RECT 2.2500 0.1575 2.3250 0.2325 ;
        RECT 1.9875 0.5175 2.0625 0.5925 ;
        RECT 1.6125 0.5100 1.6875 0.5850 ;
        RECT 1.3425 0.5850 1.4175 0.6600 ;
        RECT 1.3425 0.8100 1.4175 0.8850 ;
        RECT 1.2375 0.1800 1.3125 0.2550 ;
        RECT 1.0275 0.5100 1.1025 0.5850 ;
        RECT 0.2700 0.7125 0.3450 0.7875 ;
        LAYER M2 ;
        RECT 3.8325 0.4125 4.0875 0.4875 ;
        RECT 3.7575 0.1125 3.8325 0.4875 ;
        RECT 3.0075 0.1125 3.7575 0.1875 ;
        RECT 2.9325 0.1125 3.0075 0.7350 ;
        RECT 2.6325 0.6600 2.9325 0.7350 ;
        RECT 2.7075 0.4800 2.8575 0.5850 ;
        RECT 2.6025 0.4800 2.7075 0.5550 ;
        RECT 2.5275 0.6300 2.6325 0.7350 ;
        RECT 2.5275 0.3150 2.6025 0.5550 ;
        RECT 1.8975 0.3150 2.5275 0.3900 ;
        RECT 2.2050 0.1575 2.3700 0.2400 ;
        RECT 1.7325 0.1650 2.2050 0.2400 ;
        RECT 2.0475 0.4725 2.0775 0.6375 ;
        RECT 1.9725 0.4725 2.0475 0.8850 ;
        RECT 1.2675 0.8100 1.9725 0.8850 ;
        RECT 1.8225 0.3150 1.8975 0.7350 ;
        RECT 1.4175 0.6600 1.8225 0.7350 ;
        RECT 1.6575 0.1650 1.7325 0.5850 ;
        RECT 1.5675 0.5100 1.6575 0.5850 ;
        RECT 1.3425 0.5100 1.4175 0.7350 ;
        RECT 1.2675 0.1650 1.3575 0.2700 ;
        RECT 1.1925 0.1650 1.2675 0.8850 ;
        RECT 1.0125 0.4650 1.1175 0.7875 ;
        RECT 0.2250 0.7125 1.0125 0.7875 ;
    END
END DFSNQ_0011


MACRO DFSNQ_0111
    CLASS CORE ;
    FOREIGN DFSNQ_0111 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.8300 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN SDN
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 2.9775 0.4125 3.2925 0.4875 ;
        RECT 2.9025 0.4125 2.9775 0.9375 ;
        RECT 2.4525 0.8625 2.9025 0.9375 ;
        RECT 2.3775 0.5025 2.4525 0.9375 ;
        RECT 2.2350 0.5025 2.3775 0.6075 ;
        VIA 3.1800 0.4500 VIA12_square ;
        VIA 2.3175 0.5550 VIA12_square ;
        END
    END SDN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 4.1475 0.2925 4.4625 0.7575 ;
        VIA 4.3050 0.3525 VIA12_slot ;
        VIA 4.3050 0.6975 VIA12_slot ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.3900 0.5625 0.8550 0.6375 ;
        VIA 0.7425 0.6000 VIA12_square ;
        END
    END D
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.0375 0.4125 0.2400 0.6375 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 4.7850 -0.0750 4.8300 0.0750 ;
        RECT 4.6650 -0.0750 4.7850 0.2925 ;
        RECT 4.3650 -0.0750 4.6650 0.0750 ;
        RECT 4.2450 -0.0750 4.3650 0.2025 ;
        RECT 3.9450 -0.0750 4.2450 0.0750 ;
        RECT 3.8250 -0.0750 3.9450 0.2250 ;
        RECT 3.5025 -0.0750 3.8250 0.0750 ;
        RECT 3.4275 -0.0750 3.5025 0.2475 ;
        RECT 2.0550 -0.0750 3.4275 0.0750 ;
        RECT 1.9350 -0.0750 2.0550 0.2250 ;
        RECT 1.8450 -0.0750 1.9350 0.0750 ;
        RECT 1.7250 -0.0750 1.8450 0.2250 ;
        RECT 0.7875 -0.0750 1.7250 0.0750 ;
        RECT 0.6825 -0.0750 0.7875 0.2400 ;
        RECT 0.3750 -0.0750 0.6825 0.0750 ;
        RECT 0.2550 -0.0750 0.3750 0.1875 ;
        RECT 0.0000 -0.0750 0.2550 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 4.7850 0.9750 4.8300 1.1250 ;
        RECT 4.6650 0.6600 4.7850 1.1250 ;
        RECT 4.3650 0.9750 4.6650 1.1250 ;
        RECT 4.2450 0.8475 4.3650 1.1250 ;
        RECT 3.9450 0.9750 4.2450 1.1250 ;
        RECT 3.8250 0.8625 3.9450 1.1250 ;
        RECT 3.5250 0.9750 3.8250 1.1250 ;
        RECT 3.3975 0.8625 3.5250 1.1250 ;
        RECT 3.1050 0.9750 3.3975 1.1250 ;
        RECT 2.9850 0.8325 3.1050 1.1250 ;
        RECT 2.2650 0.9750 2.9850 1.1250 ;
        RECT 2.1450 0.8325 2.2650 1.1250 ;
        RECT 1.8450 0.9750 2.1450 1.1250 ;
        RECT 1.7250 0.8400 1.8450 1.1250 ;
        RECT 0.7875 0.9750 1.7250 1.1250 ;
        RECT 0.6825 0.8100 0.7875 1.1250 ;
        RECT 0.3750 0.9750 0.6825 1.1250 ;
        RECT 0.2550 0.8625 0.3750 1.1250 ;
        RECT 0.0000 0.9750 0.2550 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 4.6950 0.2175 4.7550 0.2775 ;
        RECT 4.6950 0.6675 4.7550 0.7275 ;
        RECT 4.6950 0.8325 4.7550 0.8925 ;
        RECT 4.5900 0.4800 4.6500 0.5400 ;
        RECT 4.4850 0.3075 4.5450 0.3675 ;
        RECT 4.4850 0.6825 4.5450 0.7425 ;
        RECT 4.3800 0.4800 4.4400 0.5400 ;
        RECT 4.2750 0.1350 4.3350 0.1950 ;
        RECT 4.2750 0.8550 4.3350 0.9150 ;
        RECT 4.1700 0.4800 4.2300 0.5400 ;
        RECT 4.0650 0.3075 4.1250 0.3675 ;
        RECT 4.0650 0.6825 4.1250 0.7425 ;
        RECT 3.9600 0.4800 4.0200 0.5400 ;
        RECT 3.8550 0.1500 3.9150 0.2100 ;
        RECT 3.8550 0.8625 3.9150 0.9225 ;
        RECT 3.7500 0.4800 3.8100 0.5400 ;
        RECT 3.6450 0.2625 3.7050 0.3225 ;
        RECT 3.6450 0.7200 3.7050 0.7800 ;
        RECT 3.5400 0.4800 3.6000 0.5400 ;
        RECT 3.4350 0.1575 3.4950 0.2175 ;
        RECT 3.4350 0.8625 3.4950 0.9225 ;
        RECT 3.3300 0.4950 3.3900 0.5550 ;
        RECT 3.2250 0.8025 3.2850 0.8625 ;
        RECT 3.1200 0.4800 3.1800 0.5400 ;
        RECT 3.0150 0.8325 3.0750 0.8925 ;
        RECT 2.9100 0.5175 2.9700 0.5775 ;
        RECT 2.8050 0.1800 2.8650 0.2400 ;
        RECT 2.8050 0.8100 2.8650 0.8700 ;
        RECT 2.7000 0.3600 2.7600 0.4200 ;
        RECT 2.5950 0.1725 2.6550 0.2325 ;
        RECT 2.5950 0.7650 2.6550 0.8250 ;
        RECT 2.4900 0.4950 2.5500 0.5550 ;
        RECT 2.3850 0.1725 2.4450 0.2325 ;
        RECT 2.3850 0.8025 2.4450 0.8625 ;
        RECT 2.2800 0.5100 2.3400 0.5700 ;
        RECT 2.1750 0.8325 2.2350 0.8925 ;
        RECT 2.0625 0.5100 2.1225 0.5700 ;
        RECT 1.9650 0.1575 2.0250 0.2175 ;
        RECT 1.9650 0.6900 2.0250 0.7500 ;
        RECT 1.8600 0.5100 1.9200 0.5700 ;
        RECT 1.7550 0.1575 1.8150 0.2175 ;
        RECT 1.7550 0.8475 1.8150 0.9075 ;
        RECT 1.6500 0.5100 1.7100 0.5700 ;
        RECT 1.4400 0.3450 1.5000 0.4050 ;
        RECT 1.4400 0.6450 1.5000 0.7050 ;
        RECT 1.3350 0.1575 1.3950 0.2175 ;
        RECT 1.3350 0.8250 1.3950 0.8850 ;
        RECT 1.2300 0.3450 1.2900 0.4050 ;
        RECT 1.1250 0.1575 1.1850 0.2175 ;
        RECT 1.1250 0.8100 1.1850 0.8700 ;
        RECT 1.0200 0.5025 1.0800 0.5625 ;
        RECT 0.9150 0.8100 0.9750 0.8700 ;
        RECT 0.8100 0.4950 0.8700 0.5550 ;
        RECT 0.7050 0.1575 0.7650 0.2175 ;
        RECT 0.7050 0.8325 0.7650 0.8925 ;
        RECT 0.4950 0.2325 0.5550 0.2925 ;
        RECT 0.4950 0.7500 0.5550 0.8100 ;
        RECT 0.3900 0.4650 0.4500 0.5250 ;
        RECT 0.2850 0.1275 0.3450 0.1875 ;
        RECT 0.2850 0.8700 0.3450 0.9300 ;
        RECT 0.1800 0.4875 0.2400 0.5475 ;
        RECT 0.0750 0.2400 0.1350 0.3000 ;
        RECT 0.0750 0.7575 0.1350 0.8175 ;
        LAYER M1 ;
        RECT 3.9675 0.4725 4.6950 0.5475 ;
        RECT 4.0575 0.2775 4.5600 0.3975 ;
        RECT 4.0575 0.6525 4.5600 0.7725 ;
        RECT 3.8925 0.3000 3.9675 0.7875 ;
        RECT 3.7125 0.3000 3.8925 0.3750 ;
        RECT 3.4575 0.7125 3.8925 0.7875 ;
        RECT 3.5325 0.4500 3.8175 0.6375 ;
        RECT 3.6375 0.2325 3.7125 0.3750 ;
        RECT 3.3825 0.4650 3.4575 0.7875 ;
        RECT 3.3300 0.4650 3.3825 0.5850 ;
        RECT 3.2025 0.6825 3.3075 0.8925 ;
        RECT 2.9175 0.1500 3.2625 0.2550 ;
        RECT 3.1050 0.3450 3.2550 0.6075 ;
        RECT 2.9100 0.6825 3.2025 0.7575 ;
        RECT 2.5950 0.4950 3.0000 0.5850 ;
        RECT 2.8050 0.1500 2.9175 0.2700 ;
        RECT 2.8050 0.6825 2.9100 0.9000 ;
        RECT 2.7375 0.3450 2.8200 0.4200 ;
        RECT 2.6700 0.3075 2.7375 0.4200 ;
        RECT 2.5200 0.6600 2.7300 0.8700 ;
        RECT 2.2050 0.1500 2.6850 0.2325 ;
        RECT 1.8000 0.3075 2.6700 0.3825 ;
        RECT 2.4900 0.4650 2.5950 0.5850 ;
        RECT 2.3400 0.6825 2.4450 0.8925 ;
        RECT 2.2050 0.4575 2.4150 0.6075 ;
        RECT 1.7250 0.6825 2.3400 0.7575 ;
        RECT 1.8000 0.4800 2.1225 0.6000 ;
        RECT 1.7250 0.3075 1.8000 0.4050 ;
        RECT 0.6000 0.3300 1.7250 0.4050 ;
        RECT 1.6500 0.4800 1.7250 0.7575 ;
        RECT 1.5750 0.4800 1.6500 0.6375 ;
        RECT 1.2900 0.8100 1.5900 0.9000 ;
        RECT 1.4175 0.6150 1.5000 0.7350 ;
        RECT 1.0800 0.1500 1.4400 0.2550 ;
        RECT 1.3425 0.4950 1.4175 0.7350 ;
        RECT 0.9825 0.4950 1.3425 0.6000 ;
        RECT 0.8925 0.7800 1.1850 0.9000 ;
        RECT 0.6825 0.4800 0.9075 0.7050 ;
        RECT 0.5250 0.2025 0.6000 0.8325 ;
        RECT 0.4725 0.2025 0.5250 0.3225 ;
        RECT 0.4725 0.7275 0.5250 0.8325 ;
        RECT 0.3900 0.4275 0.4500 0.5625 ;
        RECT 0.3150 0.2625 0.3900 0.7875 ;
        RECT 0.1425 0.2625 0.3150 0.3375 ;
        RECT 0.1650 0.7125 0.3150 0.7875 ;
        RECT 0.0675 0.7125 0.1650 0.8700 ;
        RECT 0.0675 0.2025 0.1425 0.3375 ;
        LAYER VIA1 ;
        RECT 3.6075 0.5625 3.6825 0.6375 ;
        RECT 3.0750 0.1650 3.1500 0.2400 ;
        RECT 2.5875 0.6975 2.6625 0.7725 ;
        RECT 2.5650 0.4950 2.6400 0.5700 ;
        RECT 2.2500 0.1575 2.3250 0.2325 ;
        RECT 1.9875 0.5175 2.0625 0.5925 ;
        RECT 1.6125 0.5100 1.6875 0.5850 ;
        RECT 1.3425 0.5850 1.4175 0.6600 ;
        RECT 1.3425 0.8100 1.4175 0.8850 ;
        RECT 1.2375 0.1800 1.3125 0.2550 ;
        RECT 1.0275 0.5100 1.1025 0.5850 ;
        RECT 0.2700 0.7125 0.3450 0.7875 ;
        LAYER M2 ;
        RECT 3.5175 0.5625 3.7575 0.6375 ;
        RECT 3.4425 0.1650 3.5175 0.6375 ;
        RECT 2.8275 0.1650 3.4425 0.2400 ;
        RECT 2.7525 0.1650 2.8275 0.7875 ;
        RECT 2.5275 0.6825 2.7525 0.7875 ;
        RECT 2.6025 0.4800 2.6775 0.5850 ;
        RECT 2.5275 0.3150 2.6025 0.5850 ;
        RECT 1.8975 0.3150 2.5275 0.3900 ;
        RECT 2.2050 0.1575 2.3700 0.2400 ;
        RECT 1.7325 0.1650 2.2050 0.2400 ;
        RECT 2.0475 0.4725 2.0775 0.6375 ;
        RECT 1.9725 0.4725 2.0475 0.8850 ;
        RECT 1.2675 0.8100 1.9725 0.8850 ;
        RECT 1.8225 0.3150 1.8975 0.7350 ;
        RECT 1.4175 0.6600 1.8225 0.7350 ;
        RECT 1.6575 0.1650 1.7325 0.5850 ;
        RECT 1.5675 0.5100 1.6575 0.5850 ;
        RECT 1.3425 0.5100 1.4175 0.7350 ;
        RECT 1.2675 0.1650 1.3575 0.2700 ;
        RECT 1.1925 0.1650 1.2675 0.8850 ;
        RECT 1.0125 0.4650 1.1175 0.7875 ;
        RECT 0.2250 0.7125 1.0125 0.7875 ;
    END
END DFSNQ_0111


MACRO DFSNQ_1010
    CLASS CORE ;
    FOREIGN DFSNQ_1010 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.2000 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN SDN
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 3.0825 0.4125 3.2325 0.4875 ;
        RECT 3.0075 0.4125 3.0825 0.9375 ;
        RECT 2.3325 0.8625 3.0075 0.9375 ;
        RECT 2.2575 0.4725 2.3325 0.9375 ;
        RECT 2.2275 0.4725 2.2575 0.6375 ;
        VIA 3.1200 0.4500 VIA12_square ;
        VIA 2.2800 0.5550 VIA12_square ;
        END
    END SDN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 3.5925 0.7125 3.7650 0.7875 ;
        RECT 3.5175 0.2625 3.5925 0.7875 ;
        RECT 3.0525 0.2625 3.5175 0.3375 ;
        VIA 3.6525 0.7500 VIA12_square ;
        VIA 3.5550 0.3525 VIA12_square ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.3900 0.5625 0.8550 0.6375 ;
        VIA 0.7425 0.6000 VIA12_square ;
        END
    END D
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.0375 0.4125 0.2400 0.6375 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 4.1550 -0.0750 4.2000 0.0750 ;
        RECT 4.0350 -0.0750 4.1550 0.2550 ;
        RECT 3.5250 -0.0750 4.0350 0.0750 ;
        RECT 3.4050 -0.0750 3.5250 0.2100 ;
        RECT 2.0550 -0.0750 3.4050 0.0750 ;
        RECT 1.9350 -0.0750 2.0550 0.2250 ;
        RECT 1.8450 -0.0750 1.9350 0.0750 ;
        RECT 1.7250 -0.0750 1.8450 0.2250 ;
        RECT 0.7875 -0.0750 1.7250 0.0750 ;
        RECT 0.6825 -0.0750 0.7875 0.2400 ;
        RECT 0.3750 -0.0750 0.6825 0.0750 ;
        RECT 0.2550 -0.0750 0.3750 0.1875 ;
        RECT 0.0000 -0.0750 0.2550 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 4.1550 0.9750 4.2000 1.1250 ;
        RECT 4.0500 0.6225 4.1550 1.1250 ;
        RECT 3.5250 0.9750 4.0500 1.1250 ;
        RECT 3.4050 0.8400 3.5250 1.1250 ;
        RECT 3.1050 0.9750 3.4050 1.1250 ;
        RECT 2.9850 0.8325 3.1050 1.1250 ;
        RECT 2.2650 0.9750 2.9850 1.1250 ;
        RECT 2.1450 0.8325 2.2650 1.1250 ;
        RECT 1.8450 0.9750 2.1450 1.1250 ;
        RECT 1.7250 0.8400 1.8450 1.1250 ;
        RECT 0.7875 0.9750 1.7250 1.1250 ;
        RECT 0.6825 0.8100 0.7875 1.1250 ;
        RECT 0.3750 0.9750 0.6825 1.1250 ;
        RECT 0.2550 0.8625 0.3750 1.1250 ;
        RECT 0.0000 0.9750 0.2550 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 4.0650 0.1800 4.1250 0.2400 ;
        RECT 4.0650 0.6525 4.1250 0.7125 ;
        RECT 4.0650 0.8325 4.1250 0.8925 ;
        RECT 3.9600 0.4650 4.0200 0.5250 ;
        RECT 3.8550 0.1725 3.9150 0.2325 ;
        RECT 3.8550 0.7575 3.9150 0.8175 ;
        RECT 3.6450 0.2325 3.7050 0.2925 ;
        RECT 3.6450 0.7500 3.7050 0.8100 ;
        RECT 3.5400 0.4800 3.6000 0.5400 ;
        RECT 3.4350 0.1425 3.4950 0.2025 ;
        RECT 3.4350 0.8550 3.4950 0.9150 ;
        RECT 3.3300 0.4800 3.3900 0.5400 ;
        RECT 3.2250 0.8025 3.2850 0.8625 ;
        RECT 3.1200 0.4800 3.1800 0.5400 ;
        RECT 3.0150 0.8325 3.0750 0.8925 ;
        RECT 2.9025 0.5175 2.9625 0.5775 ;
        RECT 2.8050 0.1575 2.8650 0.2175 ;
        RECT 2.8050 0.8100 2.8650 0.8700 ;
        RECT 2.7000 0.3750 2.7600 0.4350 ;
        RECT 2.5950 0.1725 2.6550 0.2325 ;
        RECT 2.5950 0.7800 2.6550 0.8400 ;
        RECT 2.4975 0.5100 2.5575 0.5700 ;
        RECT 2.3850 0.1575 2.4450 0.2175 ;
        RECT 2.3850 0.7800 2.4450 0.8400 ;
        RECT 2.2800 0.5100 2.3400 0.5700 ;
        RECT 2.1750 0.8325 2.2350 0.8925 ;
        RECT 2.0625 0.5100 2.1225 0.5700 ;
        RECT 1.9650 0.1575 2.0250 0.2175 ;
        RECT 1.9650 0.6900 2.0250 0.7500 ;
        RECT 1.8600 0.5100 1.9200 0.5700 ;
        RECT 1.7550 0.1575 1.8150 0.2175 ;
        RECT 1.7550 0.8475 1.8150 0.9075 ;
        RECT 1.6500 0.5100 1.7100 0.5700 ;
        RECT 1.4400 0.3450 1.5000 0.4050 ;
        RECT 1.4400 0.6450 1.5000 0.7050 ;
        RECT 1.3350 0.1575 1.3950 0.2175 ;
        RECT 1.3350 0.8250 1.3950 0.8850 ;
        RECT 1.2300 0.3450 1.2900 0.4050 ;
        RECT 1.1250 0.1575 1.1850 0.2175 ;
        RECT 1.1250 0.8100 1.1850 0.8700 ;
        RECT 1.0200 0.5025 1.0800 0.5625 ;
        RECT 0.9150 0.8100 0.9750 0.8700 ;
        RECT 0.8100 0.4950 0.8700 0.5550 ;
        RECT 0.7050 0.1575 0.7650 0.2175 ;
        RECT 0.7050 0.8325 0.7650 0.8925 ;
        RECT 0.4950 0.2325 0.5550 0.2925 ;
        RECT 0.4950 0.7500 0.5550 0.8100 ;
        RECT 0.3900 0.4650 0.4500 0.5250 ;
        RECT 0.2850 0.1275 0.3450 0.1875 ;
        RECT 0.2850 0.8700 0.3450 0.9300 ;
        RECT 0.1800 0.4875 0.2400 0.5475 ;
        RECT 0.0750 0.2400 0.1350 0.3000 ;
        RECT 0.0750 0.7575 0.1350 0.8175 ;
        LAYER M1 ;
        RECT 3.9300 0.3300 4.1025 0.5475 ;
        RECT 3.8550 0.7500 3.9450 0.8250 ;
        RECT 3.8550 0.1500 3.9375 0.2550 ;
        RECT 3.7800 0.1500 3.8550 0.8250 ;
        RECT 3.3000 0.4725 3.7800 0.5475 ;
        RECT 3.6000 0.1800 3.7050 0.3975 ;
        RECT 3.6000 0.6600 3.7050 0.9000 ;
        RECT 3.4575 0.3000 3.6000 0.3975 ;
        RECT 3.5100 0.6600 3.6000 0.7650 ;
        RECT 3.1875 0.6825 3.2925 0.8925 ;
        RECT 3.0375 0.3900 3.1950 0.6075 ;
        RECT 2.9100 0.6825 3.1875 0.7575 ;
        RECT 2.7600 0.1500 3.1200 0.2550 ;
        RECT 2.8500 0.4875 2.9625 0.6075 ;
        RECT 2.8050 0.6825 2.9100 0.9000 ;
        RECT 2.6025 0.5100 2.8500 0.5850 ;
        RECT 2.6700 0.3300 2.7900 0.4350 ;
        RECT 2.5800 0.6750 2.7300 0.8850 ;
        RECT 2.5650 0.1500 2.6850 0.2550 ;
        RECT 2.4975 0.3300 2.6700 0.4050 ;
        RECT 2.4975 0.4800 2.6025 0.6000 ;
        RECT 2.2800 0.1500 2.5650 0.2325 ;
        RECT 2.4225 0.3075 2.4975 0.4050 ;
        RECT 2.3775 0.6825 2.4525 0.8700 ;
        RECT 1.8000 0.3075 2.4225 0.3825 ;
        RECT 2.3325 0.4800 2.4225 0.6075 ;
        RECT 1.7250 0.6825 2.3775 0.7575 ;
        RECT 2.1975 0.4575 2.3325 0.6075 ;
        RECT 1.8000 0.4800 2.1225 0.6000 ;
        RECT 1.7250 0.3075 1.8000 0.4050 ;
        RECT 0.6000 0.3300 1.7250 0.4050 ;
        RECT 1.6500 0.4800 1.7250 0.7575 ;
        RECT 1.5750 0.4800 1.6500 0.6375 ;
        RECT 1.2900 0.8100 1.5900 0.9000 ;
        RECT 1.4175 0.6150 1.5000 0.7350 ;
        RECT 1.0800 0.1500 1.4400 0.2550 ;
        RECT 1.3425 0.4950 1.4175 0.7350 ;
        RECT 0.9825 0.4950 1.3425 0.6000 ;
        RECT 0.8925 0.7800 1.1850 0.9000 ;
        RECT 0.6825 0.4800 0.9075 0.7050 ;
        RECT 0.5250 0.2025 0.6000 0.8325 ;
        RECT 0.4725 0.2025 0.5250 0.3225 ;
        RECT 0.4725 0.7275 0.5250 0.8325 ;
        RECT 0.3900 0.4275 0.4500 0.5625 ;
        RECT 0.3150 0.2625 0.3900 0.7875 ;
        RECT 0.1425 0.2625 0.3150 0.3375 ;
        RECT 0.1650 0.7125 0.3150 0.7875 ;
        RECT 0.0675 0.7125 0.1650 0.8700 ;
        RECT 0.0675 0.2025 0.1425 0.3375 ;
        LAYER VIA1 ;
        RECT 3.9525 0.4125 4.0275 0.4875 ;
        RECT 2.8575 0.1650 2.9325 0.2400 ;
        RECT 2.6175 0.7125 2.6925 0.7875 ;
        RECT 2.5425 0.5100 2.6175 0.5850 ;
        RECT 2.3850 0.1575 2.4600 0.2325 ;
        RECT 1.9875 0.5175 2.0625 0.5925 ;
        RECT 1.6125 0.5100 1.6875 0.5850 ;
        RECT 1.3425 0.5850 1.4175 0.6600 ;
        RECT 1.3425 0.8100 1.4175 0.8850 ;
        RECT 1.2375 0.1800 1.3125 0.2550 ;
        RECT 1.0275 0.5100 1.1025 0.5850 ;
        RECT 0.2700 0.7125 0.3450 0.7875 ;
        LAYER M2 ;
        RECT 3.7425 0.4125 4.1025 0.4875 ;
        RECT 3.6675 0.1125 3.7425 0.4875 ;
        RECT 2.9325 0.1125 3.6675 0.1875 ;
        RECT 2.8575 0.1125 2.9325 0.7875 ;
        RECT 2.5725 0.7125 2.8575 0.7875 ;
        RECT 2.5425 0.5100 2.6700 0.5850 ;
        RECT 2.4675 0.3075 2.5425 0.5850 ;
        RECT 1.7325 0.1575 2.5350 0.2325 ;
        RECT 1.8975 0.3075 2.4675 0.3825 ;
        RECT 2.0475 0.4725 2.0775 0.6375 ;
        RECT 1.9725 0.4725 2.0475 0.8850 ;
        RECT 1.2675 0.8100 1.9725 0.8850 ;
        RECT 1.8225 0.3075 1.8975 0.7350 ;
        RECT 1.4175 0.6600 1.8225 0.7350 ;
        RECT 1.6575 0.1575 1.7325 0.5850 ;
        RECT 1.5675 0.5100 1.6575 0.5850 ;
        RECT 1.3425 0.5100 1.4175 0.7350 ;
        RECT 1.2675 0.1650 1.3575 0.2700 ;
        RECT 1.1925 0.1650 1.2675 0.8850 ;
        RECT 1.0125 0.4650 1.1175 0.7875 ;
        RECT 0.2250 0.7125 1.0125 0.7875 ;
    END
END DFSNQ_1010


MACRO DFSN_0011
    CLASS CORE ;
    FOREIGN DFSN_0011 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.6200 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN SDN
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 3.0900 0.4425 3.1650 0.6075 ;
        RECT 3.0150 0.4425 3.0900 0.9375 ;
        RECT 2.3325 0.8625 3.0150 0.9375 ;
        RECT 2.2575 0.4725 2.3325 0.9375 ;
        RECT 2.2275 0.4725 2.2575 0.6375 ;
        VIA 3.1125 0.5250 VIA12_square ;
        VIA 2.2800 0.5550 VIA12_square ;
        END
    END SDN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 3.7500 0.2625 3.8250 0.7875 ;
        RECT 3.2850 0.2625 3.7500 0.3375 ;
        RECT 3.6150 0.6825 3.7500 0.7875 ;
        VIA 3.6975 0.3000 VIA12_square ;
        VIA 3.6900 0.7350 VIA12_square ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 4.0500 0.4125 4.5150 0.4875 ;
        RECT 4.0050 0.2625 4.0500 0.4875 ;
        RECT 3.9000 0.2625 4.0050 0.7725 ;
        VIA 3.9750 0.3150 VIA12_square ;
        VIA 3.9525 0.6975 VIA12_square ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.3900 0.5625 0.8550 0.6375 ;
        VIA 0.7425 0.6000 VIA12_square ;
        END
    END D
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.0375 0.4125 0.2400 0.6375 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 4.3650 -0.0750 4.6200 0.0750 ;
        RECT 4.2450 -0.0750 4.3650 0.1875 ;
        RECT 3.9450 -0.0750 4.2450 0.0750 ;
        RECT 3.8250 -0.0750 3.9450 0.1875 ;
        RECT 3.5100 -0.0750 3.8250 0.0750 ;
        RECT 3.4050 -0.0750 3.5100 0.2325 ;
        RECT 2.0550 -0.0750 3.4050 0.0750 ;
        RECT 1.9350 -0.0750 2.0550 0.2250 ;
        RECT 1.8450 -0.0750 1.9350 0.0750 ;
        RECT 1.7250 -0.0750 1.8450 0.2250 ;
        RECT 0.7875 -0.0750 1.7250 0.0750 ;
        RECT 0.6825 -0.0750 0.7875 0.2400 ;
        RECT 0.3750 -0.0750 0.6825 0.0750 ;
        RECT 0.2550 -0.0750 0.3750 0.1875 ;
        RECT 0.0000 -0.0750 0.2550 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 4.3650 0.9750 4.6200 1.1250 ;
        RECT 4.2600 0.8025 4.3650 1.1250 ;
        RECT 3.9150 0.9750 4.2600 1.1250 ;
        RECT 3.8100 0.8400 3.9150 1.1250 ;
        RECT 3.5250 0.9750 3.8100 1.1250 ;
        RECT 3.4200 0.8400 3.5250 1.1250 ;
        RECT 3.1050 0.9750 3.4200 1.1250 ;
        RECT 2.9850 0.8325 3.1050 1.1250 ;
        RECT 2.2650 0.9750 2.9850 1.1250 ;
        RECT 2.1450 0.8325 2.2650 1.1250 ;
        RECT 1.8450 0.9750 2.1450 1.1250 ;
        RECT 1.7250 0.8400 1.8450 1.1250 ;
        RECT 0.7875 0.9750 1.7250 1.1250 ;
        RECT 0.6825 0.8100 0.7875 1.1250 ;
        RECT 0.3750 0.9750 0.6825 1.1250 ;
        RECT 0.2550 0.8625 0.3750 1.1250 ;
        RECT 0.0000 0.9750 0.2550 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 4.4850 0.1800 4.5450 0.2400 ;
        RECT 4.4850 0.6600 4.5450 0.7200 ;
        RECT 4.3725 0.4800 4.4325 0.5400 ;
        RECT 4.2750 0.1275 4.3350 0.1875 ;
        RECT 4.2750 0.8325 4.3350 0.8925 ;
        RECT 4.1625 0.4875 4.2225 0.5475 ;
        RECT 4.0650 0.2175 4.1250 0.2775 ;
        RECT 4.0650 0.8250 4.1250 0.8850 ;
        RECT 3.9675 0.4875 4.0275 0.5475 ;
        RECT 3.8550 0.1275 3.9150 0.1875 ;
        RECT 3.8550 0.8700 3.9150 0.9300 ;
        RECT 3.7425 0.4725 3.8025 0.5325 ;
        RECT 3.6450 0.2550 3.7050 0.3150 ;
        RECT 3.6450 0.7650 3.7050 0.8250 ;
        RECT 3.5475 0.4725 3.6075 0.5325 ;
        RECT 3.4350 0.1425 3.4950 0.2025 ;
        RECT 3.4350 0.8700 3.4950 0.9300 ;
        RECT 3.3300 0.4950 3.3900 0.5550 ;
        RECT 3.2250 0.8325 3.2850 0.8925 ;
        RECT 3.1200 0.4800 3.1800 0.5400 ;
        RECT 3.0150 0.1800 3.0750 0.2400 ;
        RECT 3.0150 0.8325 3.0750 0.8925 ;
        RECT 2.9025 0.5175 2.9625 0.5775 ;
        RECT 2.8050 0.1575 2.8650 0.2175 ;
        RECT 2.8050 0.8100 2.8650 0.8700 ;
        RECT 2.7000 0.3750 2.7600 0.4350 ;
        RECT 2.5950 0.1725 2.6550 0.2325 ;
        RECT 2.5950 0.7800 2.6550 0.8400 ;
        RECT 2.4975 0.5100 2.5575 0.5700 ;
        RECT 2.3850 0.1575 2.4450 0.2175 ;
        RECT 2.3850 0.7800 2.4450 0.8400 ;
        RECT 2.2800 0.5100 2.3400 0.5700 ;
        RECT 2.1750 0.8325 2.2350 0.8925 ;
        RECT 2.0625 0.5100 2.1225 0.5700 ;
        RECT 1.9650 0.1575 2.0250 0.2175 ;
        RECT 1.9650 0.6900 2.0250 0.7500 ;
        RECT 1.8600 0.5100 1.9200 0.5700 ;
        RECT 1.7550 0.1575 1.8150 0.2175 ;
        RECT 1.7550 0.8475 1.8150 0.9075 ;
        RECT 1.6500 0.5100 1.7100 0.5700 ;
        RECT 1.4400 0.3450 1.5000 0.4050 ;
        RECT 1.4400 0.6450 1.5000 0.7050 ;
        RECT 1.3350 0.1575 1.3950 0.2175 ;
        RECT 1.3350 0.8250 1.3950 0.8850 ;
        RECT 1.2300 0.3450 1.2900 0.4050 ;
        RECT 1.1250 0.1575 1.1850 0.2175 ;
        RECT 1.1250 0.8100 1.1850 0.8700 ;
        RECT 1.0200 0.5025 1.0800 0.5625 ;
        RECT 0.9150 0.8100 0.9750 0.8700 ;
        RECT 0.8100 0.4950 0.8700 0.5550 ;
        RECT 0.7050 0.1575 0.7650 0.2175 ;
        RECT 0.7050 0.8325 0.7650 0.8925 ;
        RECT 0.4950 0.2325 0.5550 0.2925 ;
        RECT 0.4950 0.7500 0.5550 0.8100 ;
        RECT 0.3900 0.4650 0.4500 0.5250 ;
        RECT 0.2850 0.1275 0.3450 0.1875 ;
        RECT 0.2850 0.8700 0.3450 0.9300 ;
        RECT 0.1800 0.4875 0.2400 0.5475 ;
        RECT 0.0750 0.2400 0.1350 0.3000 ;
        RECT 0.0750 0.7575 0.1350 0.8175 ;
        LAYER M1 ;
        RECT 4.5075 0.1500 4.5825 0.7275 ;
        RECT 4.4775 0.1500 4.5075 0.2700 ;
        RECT 4.2525 0.6525 4.5075 0.7275 ;
        RECT 4.4025 0.3375 4.4325 0.5700 ;
        RECT 4.3275 0.2625 4.4025 0.5700 ;
        RECT 4.2300 0.2625 4.3275 0.4050 ;
        RECT 4.1475 0.4800 4.2525 0.7275 ;
        RECT 4.0275 0.1500 4.1550 0.3675 ;
        RECT 4.0725 0.8100 4.1550 0.9000 ;
        RECT 3.9375 0.4800 4.1475 0.5550 ;
        RECT 3.9975 0.6300 4.0725 0.9000 ;
        RECT 3.8550 0.2625 4.0275 0.3675 ;
        RECT 3.8475 0.6300 3.9975 0.7650 ;
        RECT 3.5700 0.4650 3.8325 0.5475 ;
        RECT 3.6450 0.1500 3.7500 0.3900 ;
        RECT 3.6150 0.6225 3.7350 0.9000 ;
        RECT 3.5850 0.1500 3.6450 0.2550 ;
        RECT 3.4950 0.3450 3.5700 0.5475 ;
        RECT 3.4200 0.6450 3.5400 0.7500 ;
        RECT 3.3300 0.3450 3.4950 0.4200 ;
        RECT 3.3300 0.4950 3.4200 0.7500 ;
        RECT 3.2550 0.1875 3.3300 0.4200 ;
        RECT 3.3000 0.4950 3.3300 0.6000 ;
        RECT 3.2550 0.8250 3.3150 0.9000 ;
        RECT 3.1350 0.1875 3.2550 0.2700 ;
        RECT 3.1800 0.6825 3.2550 0.9000 ;
        RECT 3.0750 0.3450 3.1800 0.6075 ;
        RECT 2.9100 0.6825 3.1800 0.7575 ;
        RECT 3.0150 0.1500 3.1350 0.2700 ;
        RECT 3.0450 0.4575 3.0750 0.6075 ;
        RECT 2.9400 0.3300 2.9700 0.4125 ;
        RECT 2.8500 0.4875 2.9625 0.6075 ;
        RECT 2.8650 0.1500 2.9400 0.4125 ;
        RECT 2.8050 0.6825 2.9100 0.9000 ;
        RECT 2.7600 0.1500 2.8650 0.2550 ;
        RECT 2.6025 0.5100 2.8500 0.5850 ;
        RECT 2.6700 0.3300 2.7900 0.4350 ;
        RECT 2.5800 0.6750 2.7300 0.8850 ;
        RECT 2.5650 0.1500 2.6850 0.2550 ;
        RECT 2.4975 0.3300 2.6700 0.4050 ;
        RECT 2.4975 0.4800 2.6025 0.6000 ;
        RECT 2.2800 0.1500 2.5650 0.2325 ;
        RECT 2.4225 0.3075 2.4975 0.4050 ;
        RECT 2.3775 0.6825 2.4525 0.8700 ;
        RECT 1.8000 0.3075 2.4225 0.3825 ;
        RECT 2.3325 0.4800 2.4225 0.6075 ;
        RECT 1.7250 0.6825 2.3775 0.7575 ;
        RECT 2.1975 0.4575 2.3325 0.6075 ;
        RECT 1.8000 0.4800 2.1225 0.6000 ;
        RECT 1.7250 0.3075 1.8000 0.4050 ;
        RECT 0.6000 0.3300 1.7250 0.4050 ;
        RECT 1.6500 0.4800 1.7250 0.7575 ;
        RECT 1.5750 0.4800 1.6500 0.6375 ;
        RECT 1.2900 0.8100 1.5900 0.9000 ;
        RECT 1.4175 0.6150 1.5000 0.7350 ;
        RECT 1.0800 0.1500 1.4400 0.2550 ;
        RECT 1.3425 0.4950 1.4175 0.7350 ;
        RECT 0.9825 0.4950 1.3425 0.6000 ;
        RECT 0.8925 0.7800 1.1850 0.9000 ;
        RECT 0.6825 0.4800 0.9075 0.7050 ;
        RECT 0.5250 0.2025 0.6000 0.8325 ;
        RECT 0.4725 0.2025 0.5250 0.3225 ;
        RECT 0.4725 0.7275 0.5250 0.8325 ;
        RECT 0.3900 0.4275 0.4500 0.5625 ;
        RECT 0.3150 0.2625 0.3900 0.7875 ;
        RECT 0.1425 0.2625 0.3150 0.3375 ;
        RECT 0.1650 0.7125 0.3150 0.7875 ;
        RECT 0.0675 0.7125 0.1650 0.8700 ;
        RECT 0.0675 0.2025 0.1425 0.3375 ;
        LAYER VIA1 ;
        RECT 4.2750 0.2625 4.3500 0.3375 ;
        RECT 4.1475 0.5775 4.2225 0.6525 ;
        RECT 3.4950 0.4275 3.5700 0.5025 ;
        RECT 3.4275 0.6600 3.5025 0.7350 ;
        RECT 3.1800 0.7425 3.2550 0.8175 ;
        RECT 2.8650 0.2550 2.9400 0.3300 ;
        RECT 2.6175 0.7125 2.6925 0.7875 ;
        RECT 2.5425 0.5100 2.6175 0.5850 ;
        RECT 2.3850 0.1575 2.4600 0.2325 ;
        RECT 1.9875 0.5175 2.0625 0.5925 ;
        RECT 1.6125 0.5100 1.6875 0.5850 ;
        RECT 1.3425 0.5850 1.4175 0.6600 ;
        RECT 1.3425 0.8100 1.4175 0.8850 ;
        RECT 1.2375 0.1800 1.3125 0.2550 ;
        RECT 1.0275 0.5100 1.1025 0.5850 ;
        RECT 0.2700 0.7125 0.3450 0.7875 ;
        LAYER M2 ;
        RECT 4.2000 0.2625 4.4250 0.3375 ;
        RECT 4.1550 0.5625 4.2600 0.6675 ;
        RECT 4.1250 0.1125 4.2000 0.3375 ;
        RECT 4.0800 0.5625 4.1550 0.9375 ;
        RECT 2.9400 0.1125 4.1250 0.1875 ;
        RECT 3.5250 0.8625 4.0800 0.9375 ;
        RECT 3.4575 0.4125 3.6075 0.5325 ;
        RECT 3.4500 0.6225 3.5250 0.9375 ;
        RECT 3.3150 0.4575 3.4575 0.5325 ;
        RECT 3.4125 0.6225 3.4500 0.7725 ;
        RECT 3.2400 0.4575 3.3150 0.8550 ;
        RECT 3.1650 0.7050 3.2400 0.8550 ;
        RECT 2.8650 0.1125 2.9400 0.7875 ;
        RECT 2.5725 0.7125 2.8650 0.7875 ;
        RECT 2.5425 0.5100 2.6700 0.5850 ;
        RECT 2.4675 0.3075 2.5425 0.5850 ;
        RECT 1.7325 0.1575 2.5350 0.2325 ;
        RECT 1.8975 0.3075 2.4675 0.3825 ;
        RECT 2.0475 0.4725 2.0775 0.6375 ;
        RECT 1.9725 0.4725 2.0475 0.8850 ;
        RECT 1.2675 0.8100 1.9725 0.8850 ;
        RECT 1.8225 0.3075 1.8975 0.7350 ;
        RECT 1.4175 0.6600 1.8225 0.7350 ;
        RECT 1.6575 0.1575 1.7325 0.5850 ;
        RECT 1.5675 0.5100 1.6575 0.5850 ;
        RECT 1.3425 0.5100 1.4175 0.7350 ;
        RECT 1.2675 0.1650 1.3575 0.2700 ;
        RECT 1.1925 0.1650 1.2675 0.8850 ;
        RECT 1.0125 0.4650 1.1175 0.7875 ;
        RECT 0.2250 0.7125 1.0125 0.7875 ;
    END
END DFSN_0011


MACRO DFSN_0111
    CLASS CORE ;
    FOREIGN DFSN_0111 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.6700 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN SDN
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 3.1200 0.4800 3.2625 0.5550 ;
        RECT 3.0450 0.4800 3.1200 0.9375 ;
        RECT 2.3325 0.8625 3.0450 0.9375 ;
        RECT 2.2575 0.4725 2.3325 0.9375 ;
        RECT 2.2275 0.4725 2.2575 0.6375 ;
        VIA 3.1800 0.5175 VIA12_square ;
        VIA 2.2800 0.5550 VIA12_square ;
        END
    END SDN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 4.9875 0.2400 5.3025 0.7650 ;
        VIA 5.1450 0.3225 VIA12_slot ;
        VIA 5.1450 0.6825 VIA12_slot ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 4.1475 0.2325 4.4625 0.7350 ;
        VIA 4.3050 0.3150 VIA12_slot ;
        VIA 4.3050 0.6525 VIA12_slot ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.3900 0.5625 0.8550 0.6375 ;
        VIA 0.7425 0.6000 VIA12_square ;
        END
    END D
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.0375 0.4125 0.2400 0.6375 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 5.6025 -0.0750 5.6700 0.0750 ;
        RECT 5.5275 -0.0750 5.6025 0.3225 ;
        RECT 5.2050 -0.0750 5.5275 0.0750 ;
        RECT 5.0850 -0.0750 5.2050 0.1950 ;
        RECT 4.7700 -0.0750 5.0850 0.0750 ;
        RECT 4.6950 -0.0750 4.7700 0.2850 ;
        RECT 4.3650 -0.0750 4.6950 0.0750 ;
        RECT 4.2450 -0.0750 4.3650 0.1875 ;
        RECT 3.9450 -0.0750 4.2450 0.0750 ;
        RECT 3.8250 -0.0750 3.9450 0.2175 ;
        RECT 3.5100 -0.0750 3.8250 0.0750 ;
        RECT 3.4200 -0.0750 3.5100 0.3000 ;
        RECT 2.0550 -0.0750 3.4200 0.0750 ;
        RECT 1.9350 -0.0750 2.0550 0.2250 ;
        RECT 1.8450 -0.0750 1.9350 0.0750 ;
        RECT 1.7250 -0.0750 1.8450 0.2250 ;
        RECT 0.7875 -0.0750 1.7250 0.0750 ;
        RECT 0.6825 -0.0750 0.7875 0.2400 ;
        RECT 0.3750 -0.0750 0.6825 0.0750 ;
        RECT 0.2550 -0.0750 0.3750 0.1875 ;
        RECT 0.0000 -0.0750 0.2550 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 5.6175 0.9750 5.6700 1.1250 ;
        RECT 5.5125 0.6450 5.6175 1.1250 ;
        RECT 5.2050 0.9750 5.5125 1.1250 ;
        RECT 5.0850 0.8175 5.2050 1.1250 ;
        RECT 4.7625 0.9750 5.0850 1.1250 ;
        RECT 4.6875 0.7500 4.7625 1.1250 ;
        RECT 4.3650 0.9750 4.6875 1.1250 ;
        RECT 4.2450 0.8175 4.3650 1.1250 ;
        RECT 3.9450 0.9750 4.2450 1.1250 ;
        RECT 3.8250 0.8025 3.9450 1.1250 ;
        RECT 3.5250 0.9750 3.8250 1.1250 ;
        RECT 3.4050 0.8025 3.5250 1.1250 ;
        RECT 3.1050 0.9750 3.4050 1.1250 ;
        RECT 2.9850 0.8325 3.1050 1.1250 ;
        RECT 2.2650 0.9750 2.9850 1.1250 ;
        RECT 2.1450 0.8325 2.2650 1.1250 ;
        RECT 1.8450 0.9750 2.1450 1.1250 ;
        RECT 1.7250 0.8400 1.8450 1.1250 ;
        RECT 0.7875 0.9750 1.7250 1.1250 ;
        RECT 0.6825 0.8100 0.7875 1.1250 ;
        RECT 0.3750 0.9750 0.6825 1.1250 ;
        RECT 0.2550 0.8625 0.3750 1.1250 ;
        RECT 0.0000 0.9750 0.2550 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 5.5350 0.2325 5.5950 0.2925 ;
        RECT 5.5350 0.6675 5.5950 0.7275 ;
        RECT 5.5350 0.8325 5.5950 0.8925 ;
        RECT 5.4300 0.4800 5.4900 0.5400 ;
        RECT 5.3250 0.2925 5.3850 0.3525 ;
        RECT 5.3250 0.6600 5.3850 0.7200 ;
        RECT 5.2200 0.4800 5.2800 0.5400 ;
        RECT 5.1150 0.1350 5.1750 0.1950 ;
        RECT 5.1150 0.8325 5.1750 0.8925 ;
        RECT 5.0100 0.4800 5.0700 0.5400 ;
        RECT 4.9050 0.2925 4.9650 0.3525 ;
        RECT 4.9050 0.6600 4.9650 0.7200 ;
        RECT 4.8000 0.4800 4.8600 0.5400 ;
        RECT 4.6950 0.1950 4.7550 0.2550 ;
        RECT 4.6950 0.7950 4.7550 0.8550 ;
        RECT 4.5900 0.4725 4.6500 0.5325 ;
        RECT 4.4850 0.2850 4.5450 0.3450 ;
        RECT 4.4850 0.6525 4.5450 0.7125 ;
        RECT 4.3800 0.4725 4.4400 0.5325 ;
        RECT 4.2750 0.1275 4.3350 0.1875 ;
        RECT 4.2750 0.8325 4.3350 0.8925 ;
        RECT 4.1700 0.4725 4.2300 0.5325 ;
        RECT 4.0650 0.2850 4.1250 0.3450 ;
        RECT 4.0650 0.6525 4.1250 0.7125 ;
        RECT 3.9600 0.4725 4.0200 0.5325 ;
        RECT 3.8550 0.1425 3.9150 0.2025 ;
        RECT 3.8550 0.8175 3.9150 0.8775 ;
        RECT 3.7500 0.4875 3.8100 0.5475 ;
        RECT 3.6450 0.2400 3.7050 0.3000 ;
        RECT 3.6450 0.6600 3.7050 0.7200 ;
        RECT 3.5400 0.4875 3.6000 0.5475 ;
        RECT 3.4350 0.2100 3.4950 0.2700 ;
        RECT 3.4350 0.8175 3.4950 0.8775 ;
        RECT 3.3300 0.4875 3.3900 0.5475 ;
        RECT 3.2250 0.7350 3.2850 0.7950 ;
        RECT 3.1200 0.4875 3.1800 0.5475 ;
        RECT 3.0150 0.1800 3.0750 0.2400 ;
        RECT 3.0150 0.8325 3.0750 0.8925 ;
        RECT 2.9100 0.5100 2.9700 0.5700 ;
        RECT 2.8050 0.1575 2.8650 0.2175 ;
        RECT 2.8050 0.8100 2.8650 0.8700 ;
        RECT 2.7000 0.3750 2.7600 0.4350 ;
        RECT 2.5950 0.1725 2.6550 0.2325 ;
        RECT 2.5950 0.7800 2.6550 0.8400 ;
        RECT 2.4975 0.5100 2.5575 0.5700 ;
        RECT 2.3850 0.1575 2.4450 0.2175 ;
        RECT 2.3850 0.7800 2.4450 0.8400 ;
        RECT 2.2800 0.5100 2.3400 0.5700 ;
        RECT 2.1750 0.8325 2.2350 0.8925 ;
        RECT 2.0625 0.5100 2.1225 0.5700 ;
        RECT 1.9650 0.1575 2.0250 0.2175 ;
        RECT 1.9650 0.6900 2.0250 0.7500 ;
        RECT 1.8600 0.5100 1.9200 0.5700 ;
        RECT 1.7550 0.1575 1.8150 0.2175 ;
        RECT 1.7550 0.8475 1.8150 0.9075 ;
        RECT 1.6500 0.5100 1.7100 0.5700 ;
        RECT 1.4400 0.3450 1.5000 0.4050 ;
        RECT 1.4400 0.6450 1.5000 0.7050 ;
        RECT 1.3350 0.1575 1.3950 0.2175 ;
        RECT 1.3350 0.8250 1.3950 0.8850 ;
        RECT 1.2300 0.3450 1.2900 0.4050 ;
        RECT 1.1250 0.1575 1.1850 0.2175 ;
        RECT 1.1250 0.8100 1.1850 0.8700 ;
        RECT 1.0200 0.5025 1.0800 0.5625 ;
        RECT 0.9150 0.8100 0.9750 0.8700 ;
        RECT 0.8100 0.4950 0.8700 0.5550 ;
        RECT 0.7050 0.1575 0.7650 0.2175 ;
        RECT 0.7050 0.8325 0.7650 0.8925 ;
        RECT 0.4950 0.2325 0.5550 0.2925 ;
        RECT 0.4950 0.7500 0.5550 0.8100 ;
        RECT 0.3900 0.4650 0.4500 0.5250 ;
        RECT 0.2850 0.1275 0.3450 0.1875 ;
        RECT 0.2850 0.8700 0.3450 0.9300 ;
        RECT 0.1800 0.4875 0.2400 0.5475 ;
        RECT 0.0750 0.2400 0.1350 0.3000 ;
        RECT 0.0750 0.7575 0.1350 0.8175 ;
        LAYER M1 ;
        RECT 4.7550 0.4575 5.5200 0.5625 ;
        RECT 4.8750 0.2700 5.4150 0.3675 ;
        RECT 4.8825 0.6375 5.4075 0.7425 ;
        RECT 4.5600 0.4350 4.6800 0.5400 ;
        RECT 4.1475 0.2625 4.5750 0.3600 ;
        RECT 4.0425 0.6150 4.5675 0.7425 ;
        RECT 3.9600 0.4650 4.5600 0.5400 ;
        RECT 4.0350 0.2550 4.1475 0.3600 ;
        RECT 3.8850 0.2925 3.9600 0.7275 ;
        RECT 3.7125 0.2925 3.8850 0.3675 ;
        RECT 3.4650 0.6525 3.8850 0.7275 ;
        RECT 3.5400 0.4575 3.8100 0.5775 ;
        RECT 3.6375 0.2025 3.7125 0.3675 ;
        RECT 3.3900 0.4575 3.4650 0.7275 ;
        RECT 3.3300 0.4575 3.3900 0.5775 ;
        RECT 3.0150 0.1500 3.3300 0.2700 ;
        RECT 3.2025 0.6825 3.3075 0.8475 ;
        RECT 3.1125 0.3450 3.2550 0.6075 ;
        RECT 2.9100 0.6825 3.2025 0.7575 ;
        RECT 2.6025 0.5100 3.0000 0.5850 ;
        RECT 2.9400 0.3525 2.9775 0.4350 ;
        RECT 2.8650 0.1500 2.9400 0.4350 ;
        RECT 2.8050 0.6825 2.9100 0.9000 ;
        RECT 2.7600 0.1500 2.8650 0.2550 ;
        RECT 2.6700 0.3300 2.7900 0.4350 ;
        RECT 2.5800 0.6750 2.7300 0.8850 ;
        RECT 2.5650 0.1500 2.6850 0.2550 ;
        RECT 2.4975 0.3300 2.6700 0.4050 ;
        RECT 2.4975 0.4800 2.6025 0.6000 ;
        RECT 2.2800 0.1500 2.5650 0.2325 ;
        RECT 2.4225 0.3075 2.4975 0.4050 ;
        RECT 2.3775 0.6825 2.4525 0.8700 ;
        RECT 1.8000 0.3075 2.4225 0.3825 ;
        RECT 2.3325 0.4800 2.4225 0.6075 ;
        RECT 1.7250 0.6825 2.3775 0.7575 ;
        RECT 2.1975 0.4575 2.3325 0.6075 ;
        RECT 1.8000 0.4800 2.1225 0.6000 ;
        RECT 1.7250 0.3075 1.8000 0.4050 ;
        RECT 0.6000 0.3300 1.7250 0.4050 ;
        RECT 1.6500 0.4800 1.7250 0.7575 ;
        RECT 1.5750 0.4800 1.6500 0.6375 ;
        RECT 1.2900 0.8100 1.5900 0.9000 ;
        RECT 1.4175 0.6150 1.5000 0.7350 ;
        RECT 1.0800 0.1500 1.4400 0.2550 ;
        RECT 1.3425 0.4950 1.4175 0.7350 ;
        RECT 0.9825 0.4950 1.3425 0.6000 ;
        RECT 0.8925 0.7800 1.1850 0.9000 ;
        RECT 0.6825 0.4800 0.9075 0.7050 ;
        RECT 0.5250 0.2025 0.6000 0.8325 ;
        RECT 0.4725 0.2025 0.5250 0.3225 ;
        RECT 0.4725 0.7275 0.5250 0.8325 ;
        RECT 0.3900 0.4275 0.4500 0.5625 ;
        RECT 0.3150 0.2625 0.3900 0.7875 ;
        RECT 0.1425 0.2625 0.3150 0.3375 ;
        RECT 0.1650 0.7125 0.3150 0.7875 ;
        RECT 0.0675 0.7125 0.1650 0.8700 ;
        RECT 0.0675 0.2025 0.1425 0.3375 ;
        LAYER VIA1 ;
        RECT 4.8000 0.4725 4.8750 0.5475 ;
        RECT 3.6375 0.4800 3.7125 0.5550 ;
        RECT 3.2175 0.7275 3.2925 0.8025 ;
        RECT 3.1725 0.1650 3.2475 0.2400 ;
        RECT 2.8650 0.2925 2.9400 0.3675 ;
        RECT 2.6175 0.7125 2.6925 0.7875 ;
        RECT 2.5425 0.5100 2.6175 0.5850 ;
        RECT 2.3850 0.1575 2.4600 0.2325 ;
        RECT 1.9875 0.5175 2.0625 0.5925 ;
        RECT 1.6125 0.5100 1.6875 0.5850 ;
        RECT 1.3425 0.5850 1.4175 0.6600 ;
        RECT 1.3425 0.8100 1.4175 0.8850 ;
        RECT 1.2375 0.1800 1.3125 0.2550 ;
        RECT 1.0275 0.5100 1.1025 0.5850 ;
        RECT 0.2700 0.7125 0.3450 0.7875 ;
        LAYER M2 ;
        RECT 4.7625 0.4275 4.8900 0.5925 ;
        RECT 4.6875 0.4275 4.7625 0.8850 ;
        RECT 3.9225 0.8100 4.6875 0.8850 ;
        RECT 3.8475 0.1650 3.9225 0.8850 ;
        RECT 3.1125 0.1650 3.8475 0.2400 ;
        RECT 3.3075 0.8100 3.8475 0.8850 ;
        RECT 3.6375 0.3150 3.7125 0.6075 ;
        RECT 2.9775 0.3150 3.6375 0.3900 ;
        RECT 3.2025 0.6825 3.3075 0.8850 ;
        RECT 2.9025 0.2775 2.9775 0.3900 ;
        RECT 2.8275 0.2775 2.9025 0.7875 ;
        RECT 2.5425 0.7125 2.8275 0.7875 ;
        RECT 2.5425 0.4950 2.6700 0.6000 ;
        RECT 2.4675 0.3075 2.5425 0.6000 ;
        RECT 1.7325 0.1575 2.5350 0.2325 ;
        RECT 1.8975 0.3075 2.4675 0.3825 ;
        RECT 2.0475 0.4725 2.0775 0.6375 ;
        RECT 1.9725 0.4725 2.0475 0.8850 ;
        RECT 1.2675 0.8100 1.9725 0.8850 ;
        RECT 1.8225 0.3075 1.8975 0.7350 ;
        RECT 1.4175 0.6600 1.8225 0.7350 ;
        RECT 1.6575 0.1575 1.7325 0.5850 ;
        RECT 1.5675 0.5100 1.6575 0.5850 ;
        RECT 1.3425 0.5100 1.4175 0.7350 ;
        RECT 1.2675 0.1650 1.3575 0.2700 ;
        RECT 1.1925 0.1650 1.2675 0.8850 ;
        RECT 1.0125 0.4650 1.1175 0.7875 ;
        RECT 0.2250 0.7125 1.0125 0.7875 ;
    END
END DFSN_0111


MACRO DFSN_1010
    CLASS CORE ;
    FOREIGN DFSN_1010 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.4100 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN SDN
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 3.0525 0.4500 3.1275 0.9375 ;
        RECT 2.3325 0.8625 3.0525 0.9375 ;
        RECT 2.2575 0.4725 2.3325 0.9375 ;
        RECT 2.2275 0.4725 2.2575 0.6375 ;
        VIA 3.0900 0.5325 VIA12_square ;
        VIA 2.2800 0.5550 VIA12_square ;
        END
    END SDN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 4.2975 0.2175 4.3725 0.8325 ;
        RECT 4.2675 0.2175 4.2975 0.3825 ;
        RECT 4.2675 0.6675 4.2975 0.8325 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 3.5925 0.4125 4.0575 0.4875 ;
        RECT 3.5175 0.6750 3.6975 0.7500 ;
        RECT 3.5175 0.2625 3.5925 0.4875 ;
        RECT 3.4425 0.2625 3.5175 0.7500 ;
        VIA 3.5850 0.7125 VIA12_square ;
        VIA 3.5175 0.3525 VIA12_square ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.3900 0.5625 0.8550 0.6375 ;
        VIA 0.7425 0.6000 VIA12_square ;
        END
    END D
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.0375 0.4125 0.2400 0.6375 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 4.1550 -0.0750 4.4100 0.0750 ;
        RECT 4.0350 -0.0750 4.1550 0.1875 ;
        RECT 3.5250 -0.0750 4.0350 0.0750 ;
        RECT 3.4050 -0.0750 3.5250 0.2100 ;
        RECT 2.0550 -0.0750 3.4050 0.0750 ;
        RECT 1.9350 -0.0750 2.0550 0.2250 ;
        RECT 1.8450 -0.0750 1.9350 0.0750 ;
        RECT 1.7250 -0.0750 1.8450 0.2250 ;
        RECT 0.7875 -0.0750 1.7250 0.0750 ;
        RECT 0.6825 -0.0750 0.7875 0.2400 ;
        RECT 0.3750 -0.0750 0.6825 0.0750 ;
        RECT 0.2550 -0.0750 0.3750 0.1875 ;
        RECT 0.0000 -0.0750 0.2550 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 4.1550 0.9750 4.4100 1.1250 ;
        RECT 4.0500 0.8250 4.1550 1.1250 ;
        RECT 3.5250 0.9750 4.0500 1.1250 ;
        RECT 3.3975 0.8475 3.5250 1.1250 ;
        RECT 3.1050 0.9750 3.3975 1.1250 ;
        RECT 2.9850 0.8325 3.1050 1.1250 ;
        RECT 2.2650 0.9750 2.9850 1.1250 ;
        RECT 2.1450 0.8325 2.2650 1.1250 ;
        RECT 1.8450 0.9750 2.1450 1.1250 ;
        RECT 1.7250 0.8400 1.8450 1.1250 ;
        RECT 0.7875 0.9750 1.7250 1.1250 ;
        RECT 0.6825 0.8100 0.7875 1.1250 ;
        RECT 0.3750 0.9750 0.6825 1.1250 ;
        RECT 0.2550 0.8625 0.3750 1.1250 ;
        RECT 0.0000 0.9750 0.2550 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 4.2750 0.2700 4.3350 0.3300 ;
        RECT 4.2750 0.7200 4.3350 0.7800 ;
        RECT 4.1625 0.5100 4.2225 0.5700 ;
        RECT 4.0650 0.1275 4.1250 0.1875 ;
        RECT 4.0650 0.8550 4.1250 0.9150 ;
        RECT 3.9600 0.4650 4.0200 0.5250 ;
        RECT 3.8550 0.1725 3.9150 0.2325 ;
        RECT 3.8550 0.8325 3.9150 0.8925 ;
        RECT 3.6450 0.2325 3.7050 0.2925 ;
        RECT 3.6450 0.7500 3.7050 0.8100 ;
        RECT 3.5400 0.5100 3.6000 0.5700 ;
        RECT 3.4350 0.1425 3.4950 0.2025 ;
        RECT 3.4350 0.8550 3.4950 0.9150 ;
        RECT 3.3375 0.5325 3.3975 0.5925 ;
        RECT 3.2250 0.8025 3.2850 0.8625 ;
        RECT 3.1200 0.5100 3.1800 0.5700 ;
        RECT 3.0150 0.1800 3.0750 0.2400 ;
        RECT 3.0150 0.8325 3.0750 0.8925 ;
        RECT 2.9025 0.5175 2.9625 0.5775 ;
        RECT 2.8050 0.1575 2.8650 0.2175 ;
        RECT 2.8050 0.8100 2.8650 0.8700 ;
        RECT 2.7000 0.3750 2.7600 0.4350 ;
        RECT 2.5950 0.1725 2.6550 0.2325 ;
        RECT 2.5950 0.7800 2.6550 0.8400 ;
        RECT 2.4975 0.5100 2.5575 0.5700 ;
        RECT 2.3850 0.1575 2.4450 0.2175 ;
        RECT 2.3850 0.7800 2.4450 0.8400 ;
        RECT 2.2800 0.5100 2.3400 0.5700 ;
        RECT 2.1750 0.8325 2.2350 0.8925 ;
        RECT 2.0625 0.5100 2.1225 0.5700 ;
        RECT 1.9650 0.1575 2.0250 0.2175 ;
        RECT 1.9650 0.6900 2.0250 0.7500 ;
        RECT 1.8600 0.5100 1.9200 0.5700 ;
        RECT 1.7550 0.1575 1.8150 0.2175 ;
        RECT 1.7550 0.8475 1.8150 0.9075 ;
        RECT 1.6500 0.5100 1.7100 0.5700 ;
        RECT 1.4400 0.3450 1.5000 0.4050 ;
        RECT 1.4400 0.6450 1.5000 0.7050 ;
        RECT 1.3350 0.1575 1.3950 0.2175 ;
        RECT 1.3350 0.8250 1.3950 0.8850 ;
        RECT 1.2300 0.3450 1.2900 0.4050 ;
        RECT 1.1250 0.1575 1.1850 0.2175 ;
        RECT 1.1250 0.8100 1.1850 0.8700 ;
        RECT 1.0200 0.5025 1.0800 0.5625 ;
        RECT 0.9150 0.8100 0.9750 0.8700 ;
        RECT 0.8100 0.4950 0.8700 0.5550 ;
        RECT 0.7050 0.1575 0.7650 0.2175 ;
        RECT 0.7050 0.8325 0.7650 0.8925 ;
        RECT 0.4950 0.2325 0.5550 0.2925 ;
        RECT 0.4950 0.7500 0.5550 0.8100 ;
        RECT 0.3900 0.4650 0.4500 0.5250 ;
        RECT 0.2850 0.1275 0.3450 0.1875 ;
        RECT 0.2850 0.8700 0.3450 0.9300 ;
        RECT 0.1800 0.4875 0.2400 0.5475 ;
        RECT 0.0750 0.2400 0.1350 0.3000 ;
        RECT 0.0750 0.7575 0.1350 0.8175 ;
        LAYER M1 ;
        RECT 4.1925 0.4800 4.2225 0.6000 ;
        RECT 4.1175 0.4800 4.1925 0.7500 ;
        RECT 4.0425 0.2625 4.1850 0.4050 ;
        RECT 3.9300 0.6450 4.1175 0.7500 ;
        RECT 4.0200 0.2625 4.0425 0.5550 ;
        RECT 3.9375 0.3300 4.0200 0.5550 ;
        RECT 3.8550 0.8250 3.9450 0.9000 ;
        RECT 3.8550 0.1500 3.9375 0.2550 ;
        RECT 3.7800 0.1500 3.8550 0.9000 ;
        RECT 3.4425 0.5025 3.7800 0.5775 ;
        RECT 3.6000 0.1800 3.7050 0.4275 ;
        RECT 3.6000 0.6600 3.7050 0.9000 ;
        RECT 3.4425 0.2850 3.6000 0.4275 ;
        RECT 3.5100 0.6600 3.6000 0.7650 ;
        RECT 3.3375 0.5025 3.4425 0.6225 ;
        RECT 3.3075 0.2775 3.3675 0.3825 ;
        RECT 3.2025 0.1500 3.3075 0.3825 ;
        RECT 3.1875 0.6825 3.2925 0.8925 ;
        RECT 3.0375 0.4575 3.2625 0.6075 ;
        RECT 3.0150 0.1500 3.2025 0.2700 ;
        RECT 2.9100 0.6825 3.1875 0.7575 ;
        RECT 2.9400 0.3300 2.9700 0.4125 ;
        RECT 2.8500 0.4875 2.9625 0.6075 ;
        RECT 2.8650 0.1500 2.9400 0.4125 ;
        RECT 2.8050 0.6825 2.9100 0.9000 ;
        RECT 2.7600 0.1500 2.8650 0.2550 ;
        RECT 2.6025 0.5100 2.8500 0.5850 ;
        RECT 2.6700 0.3300 2.7900 0.4350 ;
        RECT 2.5800 0.6750 2.7300 0.8850 ;
        RECT 2.5650 0.1500 2.6850 0.2550 ;
        RECT 2.4975 0.3300 2.6700 0.4050 ;
        RECT 2.4975 0.4800 2.6025 0.6000 ;
        RECT 2.2800 0.1500 2.5650 0.2325 ;
        RECT 2.4225 0.3075 2.4975 0.4050 ;
        RECT 2.3775 0.6825 2.4525 0.8700 ;
        RECT 1.8000 0.3075 2.4225 0.3825 ;
        RECT 2.3325 0.4800 2.4225 0.6075 ;
        RECT 1.7250 0.6825 2.3775 0.7575 ;
        RECT 2.1975 0.4575 2.3325 0.6075 ;
        RECT 1.8000 0.4800 2.1225 0.6000 ;
        RECT 1.7250 0.3075 1.8000 0.4050 ;
        RECT 0.6000 0.3300 1.7250 0.4050 ;
        RECT 1.6500 0.4800 1.7250 0.7575 ;
        RECT 1.5750 0.4800 1.6500 0.6375 ;
        RECT 1.2900 0.8100 1.5900 0.9000 ;
        RECT 1.4175 0.6150 1.5000 0.7350 ;
        RECT 1.0800 0.1500 1.4400 0.2550 ;
        RECT 1.3425 0.4950 1.4175 0.7350 ;
        RECT 0.9825 0.4950 1.3425 0.6000 ;
        RECT 0.8925 0.7800 1.1850 0.9000 ;
        RECT 0.6825 0.4800 0.9075 0.7050 ;
        RECT 0.5250 0.2025 0.6000 0.8325 ;
        RECT 0.4725 0.2025 0.5250 0.3225 ;
        RECT 0.4725 0.7275 0.5250 0.8325 ;
        RECT 0.3900 0.4275 0.4500 0.5625 ;
        RECT 0.3150 0.2625 0.3900 0.7875 ;
        RECT 0.1425 0.2625 0.3150 0.3375 ;
        RECT 0.1650 0.7125 0.3150 0.7875 ;
        RECT 0.0675 0.7125 0.1650 0.8700 ;
        RECT 0.0675 0.2025 0.1425 0.3375 ;
        LAYER VIA1 ;
        RECT 4.0650 0.2625 4.1400 0.3375 ;
        RECT 3.9675 0.6600 4.0425 0.7350 ;
        RECT 3.2475 0.2925 3.3225 0.3675 ;
        RECT 3.2025 0.7350 3.2775 0.8100 ;
        RECT 2.8650 0.2550 2.9400 0.3300 ;
        RECT 2.6175 0.7125 2.6925 0.7875 ;
        RECT 2.5425 0.5100 2.6175 0.5850 ;
        RECT 2.3850 0.1575 2.4600 0.2325 ;
        RECT 1.9875 0.5175 2.0625 0.5925 ;
        RECT 1.6125 0.5100 1.6875 0.5850 ;
        RECT 1.3425 0.5850 1.4175 0.6600 ;
        RECT 1.3425 0.8100 1.4175 0.8850 ;
        RECT 1.2375 0.1800 1.3125 0.2550 ;
        RECT 1.0275 0.5100 1.1025 0.5850 ;
        RECT 0.2700 0.7125 0.3450 0.7875 ;
        LAYER M2 ;
        RECT 3.7425 0.2625 4.1850 0.3375 ;
        RECT 3.9525 0.6150 4.0575 0.9375 ;
        RECT 3.2775 0.8625 3.9525 0.9375 ;
        RECT 3.6675 0.1125 3.7425 0.3375 ;
        RECT 2.9400 0.1125 3.6675 0.1875 ;
        RECT 3.2775 0.2775 3.3675 0.3825 ;
        RECT 3.2025 0.2775 3.2775 0.9375 ;
        RECT 2.8650 0.1125 2.9400 0.7875 ;
        RECT 2.5725 0.7125 2.8650 0.7875 ;
        RECT 2.5425 0.5100 2.6700 0.5850 ;
        RECT 2.4675 0.3075 2.5425 0.5850 ;
        RECT 1.7325 0.1575 2.5350 0.2325 ;
        RECT 1.8975 0.3075 2.4675 0.3825 ;
        RECT 2.0475 0.4725 2.0775 0.6375 ;
        RECT 1.9725 0.4725 2.0475 0.8850 ;
        RECT 1.2675 0.8100 1.9725 0.8850 ;
        RECT 1.8225 0.3075 1.8975 0.7350 ;
        RECT 1.4175 0.6600 1.8225 0.7350 ;
        RECT 1.6575 0.1575 1.7325 0.5850 ;
        RECT 1.5675 0.5100 1.6575 0.5850 ;
        RECT 1.3425 0.5100 1.4175 0.7350 ;
        RECT 1.2675 0.1650 1.3575 0.2700 ;
        RECT 1.1925 0.1650 1.2675 0.8850 ;
        RECT 1.0125 0.4650 1.1175 0.7875 ;
        RECT 0.2250 0.7125 1.0125 0.7875 ;
    END
END DFSN_1010


MACRO FA1_0001
    CLASS CORE ;
    FOREIGN FA1_0001 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.2000 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 4.0875 0.1500 4.1625 0.9000 ;
        RECT 4.0575 0.1500 4.0875 0.2775 ;
        RECT 4.0350 0.8100 4.0875 0.9000 ;
        END
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 3.5925 0.7275 3.6975 0.9375 ;
        RECT 3.1575 0.8625 3.5925 0.9375 ;
        VIA 3.6450 0.8175 VIA12_square ;
        END
    END CO
    PIN CI
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 2.5875 0.3750 2.6925 0.5700 ;
        RECT 2.0325 0.4950 2.5875 0.5700 ;
        RECT 1.9575 0.4125 2.0325 0.5700 ;
        RECT 1.6050 0.4125 1.9575 0.4875 ;
        RECT 1.4400 0.4125 1.6050 0.5475 ;
        VIA 2.6400 0.4575 VIA12_square ;
        VIA 1.5225 0.4950 VIA12_square ;
        END
    END CI
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 2.2125 0.3150 2.3100 0.4200 ;
        RECT 2.1375 0.2625 2.2125 0.4200 ;
        RECT 0.9975 0.2625 2.1375 0.3375 ;
        RECT 0.8925 0.2625 0.9975 0.5475 ;
        VIA 2.2200 0.3675 VIA12_square ;
        VIA 0.9450 0.4650 VIA12_square ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 2.8425 0.5100 3.1650 0.6150 ;
        RECT 2.7675 0.5100 2.8425 0.7200 ;
        RECT 1.2825 0.6450 2.7675 0.7200 ;
        RECT 1.1775 0.4575 1.2825 0.7875 ;
        RECT 0.4650 0.7125 1.1775 0.7875 ;
        RECT 0.3900 0.4125 0.4650 0.7875 ;
        RECT 0.2850 0.4125 0.3900 0.4875 ;
        VIA 3.0825 0.5625 VIA12_square ;
        VIA 2.1450 0.6825 VIA12_square ;
        VIA 1.2300 0.5400 VIA12_square ;
        VIA 0.3675 0.4500 VIA12_square ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 3.9525 -0.0750 4.2000 0.0750 ;
        RECT 3.8175 -0.0750 3.9525 0.1875 ;
        RECT 3.1050 -0.0750 3.8175 0.0750 ;
        RECT 2.9850 -0.0750 3.1050 0.1800 ;
        RECT 2.6700 -0.0750 2.9850 0.0750 ;
        RECT 2.5950 -0.0750 2.6700 0.2100 ;
        RECT 1.0050 -0.0750 2.5950 0.0750 ;
        RECT 0.8850 -0.0750 1.0050 0.1800 ;
        RECT 0.5850 -0.0750 0.8850 0.0750 ;
        RECT 0.4650 -0.0750 0.5850 0.1800 ;
        RECT 0.1575 -0.0750 0.4650 0.0750 ;
        RECT 0.0525 -0.0750 0.1575 0.3150 ;
        RECT 0.0000 -0.0750 0.0525 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 3.9225 0.9750 4.2000 1.1250 ;
        RECT 3.8475 0.8325 3.9225 1.1250 ;
        RECT 3.1050 0.9750 3.8475 1.1250 ;
        RECT 2.9850 0.8700 3.1050 1.1250 ;
        RECT 2.6850 0.9750 2.9850 1.1250 ;
        RECT 2.5650 0.8175 2.6850 1.1250 ;
        RECT 0.9975 0.9750 2.5650 1.1250 ;
        RECT 0.8925 0.8250 0.9975 1.1250 ;
        RECT 0.5775 0.9750 0.8925 1.1250 ;
        RECT 0.4725 0.8250 0.5775 1.1250 ;
        RECT 0.1425 0.9750 0.4725 1.1250 ;
        RECT 0.0675 0.8025 0.1425 1.1250 ;
        RECT 0.0000 0.9750 0.0675 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 4.0650 0.1800 4.1250 0.2400 ;
        RECT 4.0650 0.8175 4.1250 0.8775 ;
        RECT 3.9525 0.4800 4.0125 0.5400 ;
        RECT 3.8550 0.1275 3.9150 0.1875 ;
        RECT 3.8550 0.8625 3.9150 0.9225 ;
        RECT 3.7575 0.4950 3.8175 0.5550 ;
        RECT 3.6450 0.1875 3.7050 0.2475 ;
        RECT 3.6450 0.8325 3.7050 0.8925 ;
        RECT 3.4350 0.1875 3.4950 0.2475 ;
        RECT 3.4350 0.7650 3.4950 0.8250 ;
        RECT 3.3225 0.5250 3.3825 0.5850 ;
        RECT 3.2250 0.2100 3.2850 0.2700 ;
        RECT 3.2250 0.7500 3.2850 0.8100 ;
        RECT 3.1125 0.4425 3.1725 0.5025 ;
        RECT 3.0150 0.1200 3.0750 0.1800 ;
        RECT 3.0150 0.8700 3.0750 0.9300 ;
        RECT 2.9025 0.5250 2.9625 0.5850 ;
        RECT 2.8050 0.1650 2.8650 0.2250 ;
        RECT 2.8050 0.7500 2.8650 0.8100 ;
        RECT 2.6925 0.4200 2.7525 0.4800 ;
        RECT 2.5950 0.1200 2.6550 0.1800 ;
        RECT 2.5950 0.8475 2.6550 0.9075 ;
        RECT 2.4975 0.4200 2.5575 0.4800 ;
        RECT 2.2725 0.5100 2.3325 0.5700 ;
        RECT 2.0775 0.5550 2.1375 0.6150 ;
        RECT 1.9650 0.1650 2.0250 0.2250 ;
        RECT 1.9650 0.7950 2.0250 0.8550 ;
        RECT 1.7550 0.3000 1.8150 0.3600 ;
        RECT 1.7550 0.7350 1.8150 0.7950 ;
        RECT 1.6425 0.4800 1.7025 0.5400 ;
        RECT 1.5450 0.1575 1.6050 0.2175 ;
        RECT 1.5450 0.6825 1.6050 0.7425 ;
        RECT 1.4400 0.4800 1.5000 0.5400 ;
        RECT 1.3350 0.3000 1.3950 0.3600 ;
        RECT 1.3350 0.8325 1.3950 0.8925 ;
        RECT 1.2300 0.4950 1.2900 0.5550 ;
        RECT 1.0200 0.4725 1.0800 0.5325 ;
        RECT 0.9150 0.1200 0.9750 0.1800 ;
        RECT 0.9150 0.8475 0.9750 0.9075 ;
        RECT 0.8100 0.4725 0.8700 0.5325 ;
        RECT 0.7050 0.2550 0.7650 0.3150 ;
        RECT 0.7050 0.7575 0.7650 0.8175 ;
        RECT 0.6000 0.4725 0.6600 0.5325 ;
        RECT 0.4950 0.1200 0.5550 0.1800 ;
        RECT 0.4950 0.8475 0.5550 0.9075 ;
        RECT 0.3900 0.4800 0.4500 0.5400 ;
        RECT 0.2850 0.2550 0.3450 0.3150 ;
        RECT 0.2850 0.7575 0.3450 0.8175 ;
        RECT 0.1800 0.4800 0.2400 0.5400 ;
        RECT 0.0750 0.2325 0.1350 0.2925 ;
        RECT 0.0750 0.8325 0.1350 0.8925 ;
        LAYER M1 ;
        RECT 3.9225 0.3525 4.0125 0.7050 ;
        RECT 3.7725 0.3525 3.8475 0.7275 ;
        RECT 3.7575 0.3525 3.7725 0.6225 ;
        RECT 3.6825 0.8250 3.7350 0.9000 ;
        RECT 3.6825 0.1500 3.7125 0.2775 ;
        RECT 3.6075 0.1500 3.6825 0.9000 ;
        RECT 3.4575 0.1500 3.5325 0.9000 ;
        RECT 3.4050 0.1500 3.4575 0.3150 ;
        RECT 3.4275 0.7200 3.4575 0.9000 ;
        RECT 3.2475 0.4050 3.3825 0.6450 ;
        RECT 3.2175 0.7200 3.2925 0.8400 ;
        RECT 3.2100 0.1800 3.2850 0.3300 ;
        RECT 2.8725 0.7200 3.2175 0.7950 ;
        RECT 2.8950 0.2550 3.2100 0.3300 ;
        RECT 3.0375 0.4050 3.1725 0.6450 ;
        RECT 2.8875 0.4950 2.9625 0.6450 ;
        RECT 2.7750 0.1500 2.8950 0.3300 ;
        RECT 2.3325 0.5700 2.8875 0.6450 ;
        RECT 2.7975 0.7200 2.8725 0.8400 ;
        RECT 2.6925 0.4050 2.7825 0.4950 ;
        RECT 2.4375 0.3900 2.6925 0.4950 ;
        RECT 2.4150 0.1500 2.5200 0.3150 ;
        RECT 2.0025 0.1500 2.4150 0.2250 ;
        RECT 2.2575 0.3300 2.3325 0.6450 ;
        RECT 2.1825 0.8025 2.2725 0.9000 ;
        RECT 2.1375 0.3300 2.2575 0.4050 ;
        RECT 2.1075 0.5250 2.1825 0.9000 ;
        RECT 2.0775 0.5250 2.1075 0.6450 ;
        RECT 2.0025 0.7650 2.0325 0.8850 ;
        RECT 1.9275 0.1500 2.0025 0.8850 ;
        RECT 1.7775 0.3000 1.8525 0.9000 ;
        RECT 1.3050 0.3000 1.7775 0.3750 ;
        RECT 1.7475 0.6975 1.7775 0.9000 ;
        RECT 1.6500 0.8175 1.7475 0.9000 ;
        RECT 1.4400 0.4500 1.7025 0.5850 ;
        RECT 1.3050 0.8250 1.6500 0.9000 ;
        RECT 1.1550 0.1500 1.6350 0.2250 ;
        RECT 1.5150 0.6675 1.6350 0.7425 ;
        RECT 1.4400 0.6675 1.5150 0.7500 ;
        RECT 0.7875 0.6750 1.4400 0.7500 ;
        RECT 1.1550 0.4500 1.3650 0.6000 ;
        RECT 1.0800 0.1500 1.1550 0.3375 ;
        RECT 0.7875 0.2625 1.0800 0.3375 ;
        RECT 0.5550 0.4275 1.0800 0.5700 ;
        RECT 0.6825 0.2100 0.7875 0.3375 ;
        RECT 0.6825 0.6750 0.7875 0.8400 ;
        RECT 0.3675 0.2625 0.6825 0.3375 ;
        RECT 0.3675 0.6750 0.6825 0.7500 ;
        RECT 0.1575 0.4125 0.4500 0.5850 ;
        RECT 0.2625 0.2100 0.3675 0.3375 ;
        RECT 0.2625 0.6750 0.3675 0.8400 ;
        LAYER VIA1 ;
        RECT 3.9225 0.4125 3.9975 0.4875 ;
        RECT 3.7725 0.6075 3.8475 0.6825 ;
        RECT 3.4425 0.1950 3.5175 0.2700 ;
        RECT 3.2775 0.4725 3.3525 0.5475 ;
        RECT 2.4300 0.1950 2.5050 0.2700 ;
        RECT 1.7325 0.8175 1.8075 0.8925 ;
        LAYER M2 ;
        RECT 3.5175 0.4125 4.0425 0.4875 ;
        RECT 3.7725 0.5625 3.8475 0.8100 ;
        RECT 3.3525 0.5625 3.7725 0.6375 ;
        RECT 3.4425 0.1425 3.5175 0.4875 ;
        RECT 2.5200 0.1425 3.4425 0.2175 ;
        RECT 3.2775 0.3975 3.3525 0.7875 ;
        RECT 3.0000 0.7125 3.2775 0.7875 ;
        RECT 2.9250 0.7125 3.0000 0.9375 ;
        RECT 1.8525 0.8625 2.9250 0.9375 ;
        RECT 2.4150 0.1425 2.5200 0.3150 ;
        RECT 1.6875 0.8025 1.8525 0.9375 ;
    END
END FA1_0001


MACRO FA1_0011
    CLASS CORE ;
    FOREIGN FA1_0011 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.9900 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 3.8775 0.3075 3.9525 0.7425 ;
        RECT 3.7125 0.3075 3.8775 0.3825 ;
        RECT 3.7125 0.6675 3.8775 0.7425 ;
        RECT 3.6375 0.2175 3.7125 0.3825 ;
        RECT 3.6375 0.6675 3.7125 0.8325 ;
        END
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 3.2475 0.2625 3.3225 0.9375 ;
        RECT 3.1125 0.2625 3.2475 0.3375 ;
        RECT 2.4900 0.8625 3.2475 0.9375 ;
        VIA 3.2850 0.7725 VIA12_square ;
        VIA 3.1950 0.3000 VIA12_square ;
        END
    END CO
    PIN CI
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.9425 0.3750 2.0475 0.5925 ;
        RECT 1.5150 0.5175 1.9425 0.5925 ;
        RECT 1.4400 0.2625 1.5150 0.5925 ;
        RECT 1.2300 0.2625 1.4400 0.3375 ;
        RECT 1.0800 0.2625 1.2300 0.4350 ;
        RECT 0.8250 0.2625 1.0800 0.3375 ;
        VIA 1.9950 0.4575 VIA12_square ;
        VIA 1.1550 0.3825 VIA12_square ;
        END
    END CI
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.6650 0.3600 1.7625 0.4350 ;
        RECT 1.5900 0.1125 1.6650 0.4350 ;
        RECT 0.5850 0.1125 1.5900 0.1875 ;
        RECT 0.5100 0.1125 0.5850 0.4875 ;
        RECT 0.3600 0.4125 0.5100 0.4875 ;
        VIA 1.6800 0.3975 VIA12_square ;
        VIA 0.4725 0.4500 VIA12_square ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 2.3700 0.4725 2.5425 0.5775 ;
        RECT 2.2950 0.4725 2.3700 0.8925 ;
        RECT 1.5450 0.8175 2.2950 0.8925 ;
        RECT 1.4700 0.8175 1.5450 0.9375 ;
        RECT 0.9300 0.8625 1.4700 0.9375 ;
        RECT 0.8550 0.8175 0.9300 0.9375 ;
        RECT 0.7050 0.8175 0.8550 0.8925 ;
        VIA 2.4600 0.5250 VIA12_square ;
        VIA 1.5825 0.8550 VIA12_square ;
        VIA 0.8175 0.8550 VIA12_square ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 3.9450 -0.0750 3.9900 0.0750 ;
        RECT 3.8250 -0.0750 3.9450 0.2325 ;
        RECT 3.5100 -0.0750 3.8250 0.0750 ;
        RECT 3.4200 -0.0750 3.5100 0.3075 ;
        RECT 3.0825 -0.0750 3.4200 0.0750 ;
        RECT 3.0075 -0.0750 3.0825 0.3150 ;
        RECT 2.4750 -0.0750 3.0075 0.0750 ;
        RECT 2.3550 -0.0750 2.4750 0.1800 ;
        RECT 2.0325 -0.0750 2.3550 0.0750 ;
        RECT 1.9575 -0.0750 2.0325 0.2625 ;
        RECT 0.5850 -0.0750 1.9575 0.0750 ;
        RECT 0.4650 -0.0750 0.5850 0.1800 ;
        RECT 0.1425 -0.0750 0.4650 0.0750 ;
        RECT 0.0675 -0.0750 0.1425 0.3075 ;
        RECT 0.0000 -0.0750 0.0675 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 3.9450 0.9750 3.9900 1.1250 ;
        RECT 3.8250 0.8175 3.9450 1.1250 ;
        RECT 3.5175 0.9750 3.8250 1.1250 ;
        RECT 3.4125 0.6675 3.5175 1.1250 ;
        RECT 3.0975 0.9750 3.4125 1.1250 ;
        RECT 2.9925 0.6450 3.0975 1.1250 ;
        RECT 2.4750 0.9750 2.9925 1.1250 ;
        RECT 2.3550 0.8700 2.4750 1.1250 ;
        RECT 2.0550 0.9750 2.3550 1.1250 ;
        RECT 1.9350 0.8025 2.0550 1.1250 ;
        RECT 0.5625 0.9750 1.9350 1.1250 ;
        RECT 0.4875 0.7800 0.5625 1.1250 ;
        RECT 0.1425 0.9750 0.4875 1.1250 ;
        RECT 0.0675 0.7875 0.1425 1.1250 ;
        RECT 0.0000 0.9750 0.0675 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 3.8550 0.1575 3.9150 0.2175 ;
        RECT 3.8550 0.8325 3.9150 0.8925 ;
        RECT 3.7425 0.4875 3.8025 0.5475 ;
        RECT 3.6450 0.2700 3.7050 0.3300 ;
        RECT 3.6450 0.7200 3.7050 0.7800 ;
        RECT 3.5400 0.4875 3.6000 0.5475 ;
        RECT 3.4350 0.2025 3.4950 0.2625 ;
        RECT 3.4350 0.6900 3.4950 0.7500 ;
        RECT 3.4350 0.8550 3.4950 0.9150 ;
        RECT 3.3300 0.4950 3.3900 0.5550 ;
        RECT 3.2250 0.2175 3.2850 0.2775 ;
        RECT 3.2250 0.7500 3.2850 0.8100 ;
        RECT 3.1200 0.4950 3.1800 0.5550 ;
        RECT 3.0150 0.2025 3.0750 0.2625 ;
        RECT 3.0150 0.6675 3.0750 0.7275 ;
        RECT 3.0150 0.8325 3.0750 0.8925 ;
        RECT 2.8050 0.1950 2.8650 0.2550 ;
        RECT 2.8050 0.7800 2.8650 0.8400 ;
        RECT 2.7000 0.5025 2.7600 0.5625 ;
        RECT 2.5950 0.2100 2.6550 0.2700 ;
        RECT 2.5950 0.7800 2.6550 0.8400 ;
        RECT 2.4900 0.5100 2.5500 0.5700 ;
        RECT 2.3850 0.1200 2.4450 0.1800 ;
        RECT 2.3850 0.8700 2.4450 0.9300 ;
        RECT 2.2800 0.5100 2.3400 0.5700 ;
        RECT 2.1750 0.1950 2.2350 0.2550 ;
        RECT 2.1750 0.7875 2.2350 0.8475 ;
        RECT 2.0625 0.4200 2.1225 0.4800 ;
        RECT 1.9650 0.1725 2.0250 0.2325 ;
        RECT 1.9650 0.8250 2.0250 0.8850 ;
        RECT 1.8675 0.4200 1.9275 0.4800 ;
        RECT 1.6500 0.5100 1.7100 0.5700 ;
        RECT 1.4400 0.5100 1.5000 0.5700 ;
        RECT 1.3350 0.1950 1.3950 0.2550 ;
        RECT 1.3350 0.7800 1.3950 0.8400 ;
        RECT 1.1250 0.1575 1.1850 0.2175 ;
        RECT 1.1250 0.6825 1.1850 0.7425 ;
        RECT 1.0200 0.4725 1.0800 0.5325 ;
        RECT 0.9150 0.3000 0.9750 0.3600 ;
        RECT 0.9150 0.6450 0.9750 0.7050 ;
        RECT 0.8100 0.8400 0.8700 0.9000 ;
        RECT 0.6000 0.4275 0.6600 0.4875 ;
        RECT 0.4950 0.1200 0.5550 0.1800 ;
        RECT 0.4950 0.8325 0.5550 0.8925 ;
        RECT 0.3900 0.4275 0.4500 0.4875 ;
        RECT 0.2850 0.2550 0.3450 0.3150 ;
        RECT 0.2850 0.7200 0.3450 0.7800 ;
        RECT 0.1800 0.4800 0.2400 0.5400 ;
        RECT 0.0750 0.2025 0.1350 0.2625 ;
        RECT 0.0750 0.8325 0.1350 0.8925 ;
        LAYER M1 ;
        RECT 3.5475 0.4575 3.8025 0.5775 ;
        RECT 3.4725 0.4125 3.5475 0.5775 ;
        RECT 3.2850 0.4650 3.3900 0.5850 ;
        RECT 3.1800 0.6600 3.3300 0.8925 ;
        RECT 3.1575 0.1800 3.3225 0.3900 ;
        RECT 2.9100 0.4875 3.2850 0.5700 ;
        RECT 2.7375 0.4875 2.9100 0.5775 ;
        RECT 2.8125 0.1500 2.8875 0.3825 ;
        RECT 2.7375 0.6525 2.8875 0.9000 ;
        RECT 2.7300 0.1500 2.8125 0.3450 ;
        RECT 2.6325 0.4200 2.7375 0.5775 ;
        RECT 2.5725 0.7200 2.6625 0.8700 ;
        RECT 2.5800 0.1800 2.6550 0.3300 ;
        RECT 2.2575 0.2550 2.5800 0.3300 ;
        RECT 2.2575 0.7200 2.5725 0.7950 ;
        RECT 2.4225 0.4050 2.5575 0.6450 ;
        RECT 2.2725 0.4650 2.3475 0.6450 ;
        RECT 1.7175 0.5700 2.2725 0.6450 ;
        RECT 2.1525 0.1725 2.2575 0.3300 ;
        RECT 2.1525 0.7200 2.2575 0.8700 ;
        RECT 1.9425 0.4050 2.1675 0.4950 ;
        RECT 1.8225 0.4200 1.9425 0.4950 ;
        RECT 1.8075 0.1500 1.8825 0.3150 ;
        RECT 1.4025 0.1500 1.8075 0.2250 ;
        RECT 1.6425 0.3000 1.7175 0.6450 ;
        RECT 1.5525 0.7875 1.6650 0.9000 ;
        RECT 1.6125 0.3000 1.6425 0.3750 ;
        RECT 1.4775 0.4650 1.5525 0.9000 ;
        RECT 1.4400 0.4650 1.4775 0.6075 ;
        RECT 1.3650 0.1500 1.4025 0.3750 ;
        RECT 1.3650 0.6825 1.4025 0.8700 ;
        RECT 1.3275 0.1500 1.3650 0.8700 ;
        RECT 1.2900 0.3000 1.3275 0.7575 ;
        RECT 0.7350 0.1500 1.2150 0.2250 ;
        RECT 1.1100 0.3000 1.2150 0.5325 ;
        RECT 1.0500 0.6075 1.2150 0.8325 ;
        RECT 0.9900 0.4575 1.1100 0.5325 ;
        RECT 0.8850 0.3000 1.0050 0.3750 ;
        RECT 0.8850 0.6150 0.9750 0.7350 ;
        RECT 0.7350 0.8175 0.9000 0.9000 ;
        RECT 0.8100 0.3000 0.8850 0.7350 ;
        RECT 0.6600 0.1500 0.7350 0.3300 ;
        RECT 0.6600 0.5625 0.7350 0.9000 ;
        RECT 0.3450 0.4050 0.7050 0.4875 ;
        RECT 0.2550 0.2550 0.6600 0.3300 ;
        RECT 0.2400 0.5625 0.6600 0.6375 ;
        RECT 0.2175 0.7125 0.4125 0.8775 ;
        RECT 0.1650 0.4350 0.2400 0.6375 ;
        LAYER VIA1 ;
        RECT 3.4725 0.4575 3.5475 0.5325 ;
        RECT 2.7675 0.1650 2.8425 0.2400 ;
        RECT 2.7675 0.6975 2.8425 0.7725 ;
        RECT 2.6475 0.4575 2.7225 0.5325 ;
        RECT 1.8075 0.1950 1.8825 0.2700 ;
        RECT 1.0950 0.6750 1.1700 0.7500 ;
        RECT 0.8100 0.5100 0.8850 0.5850 ;
        RECT 0.2775 0.7125 0.3525 0.7875 ;
        LAYER M2 ;
        RECT 3.4725 0.1125 3.5475 0.5775 ;
        RECT 2.8875 0.1125 3.4725 0.1875 ;
        RECT 2.8125 0.1125 2.8875 0.7875 ;
        RECT 1.9275 0.1650 2.8125 0.2400 ;
        RECT 2.7300 0.6825 2.8125 0.7875 ;
        RECT 2.6325 0.3150 2.7375 0.5775 ;
        RECT 2.2050 0.3150 2.6325 0.3900 ;
        RECT 2.1300 0.3150 2.2050 0.7425 ;
        RECT 1.3650 0.6675 2.1300 0.7425 ;
        RECT 1.7625 0.1650 1.9275 0.2850 ;
        RECT 1.2900 0.5100 1.3650 0.7425 ;
        RECT 0.7350 0.5100 1.2900 0.5850 ;
        RECT 1.0500 0.6600 1.2150 0.7650 ;
        RECT 0.3675 0.6600 1.0500 0.7350 ;
        RECT 0.2625 0.6600 0.3675 0.8325 ;
    END
END FA1_0011


MACRO FA1_0111
    CLASS CORE ;
    FOREIGN FA1_0111 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.0900 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 5.4075 0.2625 5.7225 0.7275 ;
        VIA 5.5650 0.3225 VIA12_slot ;
        VIA 5.5650 0.6675 VIA12_slot ;
        END
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 4.5675 0.2625 4.8825 0.7125 ;
        VIA 4.7250 0.3225 VIA12_slot ;
        VIA 4.7250 0.6525 VIA12_slot ;
        END
    END CO
    PIN CI
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 3.2925 0.2625 3.7575 0.3375 ;
        RECT 3.2175 0.2625 3.2925 0.5775 ;
        RECT 2.4750 0.5025 3.2175 0.5775 ;
        RECT 2.3250 0.4725 2.4750 0.5775 ;
        VIA 3.2550 0.4500 VIA12_square ;
        VIA 2.4000 0.5250 VIA12_square ;
        END
    END CI
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 2.7975 0.3000 2.9400 0.4050 ;
        RECT 2.7150 0.1650 2.7975 0.4050 ;
        RECT 1.7550 0.1650 2.7150 0.2400 ;
        RECT 1.7550 0.4875 1.8450 0.5625 ;
        RECT 1.6800 0.1650 1.7550 0.5625 ;
        RECT 0.9975 0.1650 1.6800 0.2400 ;
        RECT 0.8925 0.1650 0.9975 0.5625 ;
        RECT 0.4275 0.2625 0.8925 0.3375 ;
        RECT 0.3525 0.2625 0.4275 0.4875 ;
        RECT 0.1050 0.4125 0.3525 0.4875 ;
        VIA 2.8575 0.3525 VIA12_square ;
        VIA 1.7625 0.5250 VIA12_square ;
        VIA 0.9450 0.4875 VIA12_square ;
        VIA 0.2175 0.4500 VIA12_square ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 3.7200 0.5625 3.8400 0.6375 ;
        RECT 3.6450 0.5625 3.7200 0.8775 ;
        RECT 1.1925 0.8025 3.6450 0.8775 ;
        RECT 1.1925 0.4725 1.3425 0.5775 ;
        RECT 1.1175 0.4725 1.1925 0.8775 ;
        RECT 0.6075 0.7125 1.1175 0.7875 ;
        RECT 0.5025 0.4350 0.6075 0.7875 ;
        VIA 3.7575 0.6000 VIA12_square ;
        VIA 2.8425 0.8400 VIA12_square ;
        VIA 1.2675 0.5250 VIA12_square ;
        VIA 0.5550 0.5100 VIA12_square ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 6.0225 -0.0750 6.0900 0.0750 ;
        RECT 5.9475 -0.0750 6.0225 0.3075 ;
        RECT 5.6250 -0.0750 5.9475 0.0750 ;
        RECT 5.5050 -0.0750 5.6250 0.2025 ;
        RECT 5.2050 -0.0750 5.5050 0.0750 ;
        RECT 5.0850 -0.0750 5.2050 0.3675 ;
        RECT 4.7850 -0.0750 5.0850 0.0750 ;
        RECT 4.6650 -0.0750 4.7850 0.2025 ;
        RECT 4.3425 -0.0750 4.6650 0.0750 ;
        RECT 4.2675 -0.0750 4.3425 0.3150 ;
        RECT 3.7350 -0.0750 4.2675 0.0750 ;
        RECT 3.6150 -0.0750 3.7350 0.1800 ;
        RECT 3.3000 -0.0750 3.6150 0.0750 ;
        RECT 3.2250 -0.0750 3.3000 0.2625 ;
        RECT 1.8375 -0.0750 3.2250 0.0750 ;
        RECT 1.7325 -0.0750 1.8375 0.2400 ;
        RECT 0.9975 -0.0750 1.7325 0.0750 ;
        RECT 0.8775 -0.0750 0.9975 0.2100 ;
        RECT 0.5850 -0.0750 0.8775 0.0750 ;
        RECT 0.4650 -0.0750 0.5850 0.1875 ;
        RECT 0.1425 -0.0750 0.4650 0.0750 ;
        RECT 0.0675 -0.0750 0.1425 0.3000 ;
        RECT 0.0000 -0.0750 0.0675 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 6.0225 0.9750 6.0900 1.1250 ;
        RECT 5.9475 0.6375 6.0225 1.1250 ;
        RECT 5.6175 0.9750 5.9475 1.1250 ;
        RECT 5.5125 0.7875 5.6175 1.1250 ;
        RECT 5.2050 0.9750 5.5125 1.1250 ;
        RECT 5.0850 0.6600 5.2050 1.1250 ;
        RECT 4.7775 0.9750 5.0850 1.1250 ;
        RECT 4.6725 0.7875 4.7775 1.1250 ;
        RECT 4.3650 0.9750 4.6725 1.1250 ;
        RECT 4.2450 0.6600 4.3650 1.1250 ;
        RECT 3.7350 0.9750 4.2450 1.1250 ;
        RECT 3.6150 0.8700 3.7350 1.1250 ;
        RECT 3.3150 0.9750 3.6150 1.1250 ;
        RECT 3.1950 0.8025 3.3150 1.1250 ;
        RECT 1.8600 0.9750 3.1950 1.1250 ;
        RECT 1.7325 0.8100 1.8600 1.1250 ;
        RECT 0.9975 0.9750 1.7325 1.1250 ;
        RECT 0.8850 0.8175 0.9975 1.1250 ;
        RECT 0.5850 0.9750 0.8850 1.1250 ;
        RECT 0.4650 0.8175 0.5850 1.1250 ;
        RECT 0.1575 0.9750 0.4650 1.1250 ;
        RECT 0.0525 0.6450 0.1575 1.1250 ;
        RECT 0.0000 0.9750 0.0525 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 5.9550 0.2100 6.0150 0.2700 ;
        RECT 5.9550 0.6675 6.0150 0.7275 ;
        RECT 5.9550 0.8325 6.0150 0.8925 ;
        RECT 5.8500 0.4650 5.9100 0.5250 ;
        RECT 5.7450 0.2250 5.8050 0.2850 ;
        RECT 5.7450 0.7575 5.8050 0.8175 ;
        RECT 5.6400 0.4650 5.7000 0.5250 ;
        RECT 5.5350 0.1275 5.5950 0.1875 ;
        RECT 5.5350 0.8175 5.5950 0.8775 ;
        RECT 5.4300 0.4650 5.4900 0.5250 ;
        RECT 5.3250 0.2250 5.3850 0.2850 ;
        RECT 5.3250 0.7575 5.3850 0.8175 ;
        RECT 5.2200 0.4725 5.2800 0.5325 ;
        RECT 5.1150 0.1200 5.1750 0.1800 ;
        RECT 5.1150 0.2850 5.1750 0.3450 ;
        RECT 5.1150 0.6900 5.1750 0.7500 ;
        RECT 5.1150 0.8550 5.1750 0.9150 ;
        RECT 5.0100 0.4725 5.0700 0.5325 ;
        RECT 4.9050 0.2250 4.9650 0.2850 ;
        RECT 4.9050 0.7575 4.9650 0.8175 ;
        RECT 4.8000 0.4650 4.8600 0.5250 ;
        RECT 4.6950 0.1275 4.7550 0.1875 ;
        RECT 4.6950 0.8175 4.7550 0.8775 ;
        RECT 4.5900 0.4650 4.6500 0.5250 ;
        RECT 4.4850 0.2250 4.5450 0.2850 ;
        RECT 4.4850 0.7575 4.5450 0.8175 ;
        RECT 4.3800 0.4650 4.4400 0.5250 ;
        RECT 4.2750 0.2100 4.3350 0.2700 ;
        RECT 4.2750 0.6675 4.3350 0.7275 ;
        RECT 4.2750 0.8325 4.3350 0.8925 ;
        RECT 4.0650 0.1800 4.1250 0.2400 ;
        RECT 4.0650 0.7800 4.1250 0.8400 ;
        RECT 3.9600 0.4725 4.0200 0.5325 ;
        RECT 3.8550 0.1950 3.9150 0.2550 ;
        RECT 3.8550 0.8025 3.9150 0.8625 ;
        RECT 3.7500 0.5100 3.8100 0.5700 ;
        RECT 3.6450 0.1200 3.7050 0.1800 ;
        RECT 3.6450 0.8700 3.7050 0.9300 ;
        RECT 3.5325 0.5100 3.5925 0.5700 ;
        RECT 3.4350 0.1950 3.4950 0.2550 ;
        RECT 3.4350 0.7875 3.4950 0.8475 ;
        RECT 3.3225 0.4200 3.3825 0.4800 ;
        RECT 3.2250 0.1725 3.2850 0.2325 ;
        RECT 3.2250 0.8325 3.2850 0.8925 ;
        RECT 3.1200 0.4200 3.1800 0.4800 ;
        RECT 2.9100 0.5100 2.9700 0.5700 ;
        RECT 2.7000 0.5250 2.7600 0.5850 ;
        RECT 2.5950 0.1950 2.6550 0.2550 ;
        RECT 2.5950 0.7800 2.6550 0.8400 ;
        RECT 2.3850 0.1575 2.4450 0.2175 ;
        RECT 2.3850 0.8325 2.4450 0.8925 ;
        RECT 2.2800 0.4950 2.3400 0.5550 ;
        RECT 2.1750 0.3225 2.2350 0.3825 ;
        RECT 2.1750 0.6675 2.2350 0.7275 ;
        RECT 2.0700 0.4950 2.1300 0.5550 ;
        RECT 1.9650 0.2400 2.0250 0.3000 ;
        RECT 1.9650 0.7500 2.0250 0.8100 ;
        RECT 1.7550 0.1575 1.8150 0.2175 ;
        RECT 1.7550 0.8325 1.8150 0.8925 ;
        RECT 1.6500 0.4950 1.7100 0.5550 ;
        RECT 1.4400 0.4950 1.5000 0.5550 ;
        RECT 1.3350 0.3225 1.3950 0.3825 ;
        RECT 1.3350 0.6675 1.3950 0.7275 ;
        RECT 1.2300 0.4950 1.2900 0.5550 ;
        RECT 1.0200 0.4725 1.0800 0.5325 ;
        RECT 0.9150 0.1275 0.9750 0.1875 ;
        RECT 0.9150 0.8400 0.9750 0.9000 ;
        RECT 0.8100 0.4725 0.8700 0.5325 ;
        RECT 0.7050 0.2775 0.7650 0.3375 ;
        RECT 0.7050 0.6750 0.7650 0.7350 ;
        RECT 0.6000 0.4725 0.6600 0.5325 ;
        RECT 0.4950 0.1200 0.5550 0.1800 ;
        RECT 0.4950 0.8400 0.5550 0.9000 ;
        RECT 0.3900 0.4725 0.4500 0.5325 ;
        RECT 0.2850 0.2700 0.3450 0.3300 ;
        RECT 0.2850 0.6975 0.3450 0.7575 ;
        RECT 0.1800 0.4725 0.2400 0.5325 ;
        RECT 0.0750 0.1950 0.1350 0.2550 ;
        RECT 0.0750 0.6675 0.1350 0.7275 ;
        RECT 0.0750 0.8325 0.1350 0.8925 ;
        LAYER M1 ;
        RECT 5.1750 0.4425 5.9400 0.5475 ;
        RECT 5.7225 0.1950 5.8275 0.3675 ;
        RECT 5.7375 0.6225 5.8125 0.8700 ;
        RECT 5.3925 0.6225 5.7375 0.7125 ;
        RECT 5.4075 0.2775 5.7225 0.3675 ;
        RECT 5.3025 0.1950 5.4075 0.3675 ;
        RECT 5.3175 0.6225 5.3925 0.8700 ;
        RECT 5.0250 0.4425 5.1000 0.5475 ;
        RECT 4.0575 0.4425 5.0250 0.5325 ;
        RECT 4.8825 0.1950 4.9875 0.3675 ;
        RECT 4.8975 0.6075 4.9725 0.8700 ;
        RECT 4.5525 0.6075 4.8975 0.6975 ;
        RECT 4.5675 0.2775 4.8825 0.3675 ;
        RECT 4.4625 0.1950 4.5675 0.3675 ;
        RECT 4.4775 0.6075 4.5525 0.8700 ;
        RECT 4.0275 0.1500 4.1925 0.3450 ;
        RECT 4.0200 0.6525 4.1700 0.9000 ;
        RECT 3.9525 0.4425 4.0575 0.5625 ;
        RECT 3.8325 0.1725 3.9375 0.3300 ;
        RECT 3.8325 0.7200 3.9375 0.8850 ;
        RECT 3.6675 0.4050 3.8475 0.6450 ;
        RECT 3.5175 0.2550 3.8325 0.3300 ;
        RECT 3.5175 0.7200 3.8325 0.7950 ;
        RECT 3.5175 0.4650 3.5925 0.6450 ;
        RECT 3.4125 0.1725 3.5175 0.3300 ;
        RECT 2.9700 0.5700 3.5175 0.6450 ;
        RECT 3.4125 0.7200 3.5175 0.8700 ;
        RECT 3.2625 0.4050 3.4125 0.4950 ;
        RECT 3.0525 0.3900 3.2625 0.4950 ;
        RECT 3.0450 0.1650 3.1500 0.3150 ;
        RECT 2.6625 0.1650 3.0450 0.2400 ;
        RECT 2.8950 0.3150 2.9700 0.6450 ;
        RECT 2.8200 0.7875 2.9250 0.9000 ;
        RECT 2.7675 0.3150 2.8950 0.3900 ;
        RECT 2.7375 0.4950 2.8200 0.9000 ;
        RECT 2.7000 0.4950 2.7375 0.6150 ;
        RECT 2.6250 0.1650 2.6625 0.3900 ;
        RECT 2.6250 0.6900 2.6625 0.8700 ;
        RECT 2.5875 0.1650 2.6250 0.8700 ;
        RECT 2.5500 0.3150 2.5875 0.7650 ;
        RECT 2.0325 0.1500 2.4750 0.2250 ;
        RECT 2.3100 0.4725 2.4750 0.5775 ;
        RECT 2.0325 0.8250 2.4750 0.9000 ;
        RECT 2.2725 0.3000 2.4450 0.3900 ;
        RECT 2.2725 0.6525 2.4450 0.7500 ;
        RECT 2.0400 0.4800 2.3100 0.5700 ;
        RECT 2.1075 0.3000 2.2725 0.4050 ;
        RECT 2.1075 0.6450 2.2725 0.7500 ;
        RECT 1.9575 0.1500 2.0325 0.3900 ;
        RECT 1.9575 0.6600 2.0325 0.9000 ;
        RECT 1.6575 0.3150 1.9575 0.3900 ;
        RECT 1.6575 0.6600 1.9575 0.7350 ;
        RECT 1.6500 0.4650 1.9350 0.5850 ;
        RECT 1.5825 0.1500 1.6575 0.3900 ;
        RECT 1.5825 0.6600 1.6575 0.9000 ;
        RECT 1.1475 0.1500 1.5825 0.2250 ;
        RECT 1.1475 0.8250 1.5825 0.9000 ;
        RECT 1.1850 0.4875 1.5450 0.5625 ;
        RECT 1.2225 0.3000 1.5075 0.4125 ;
        RECT 1.2225 0.6375 1.5075 0.7500 ;
        RECT 1.0725 0.1500 1.1475 0.3600 ;
        RECT 1.0725 0.6675 1.1475 0.9000 ;
        RECT 0.8025 0.4350 1.0800 0.5850 ;
        RECT 0.8025 0.2850 1.0725 0.3600 ;
        RECT 0.3600 0.6675 1.0725 0.7425 ;
        RECT 0.6675 0.2625 0.8025 0.3600 ;
        RECT 0.2475 0.2625 0.6675 0.3375 ;
        RECT 0.3900 0.4350 0.6675 0.5850 ;
        RECT 0.2700 0.6675 0.3600 0.7875 ;
        RECT 0.0675 0.4125 0.3150 0.5700 ;
        LAYER VIA1 ;
        RECT 5.2125 0.4575 5.2875 0.5325 ;
        RECT 4.0725 0.2100 4.1475 0.2850 ;
        RECT 4.0575 0.4575 4.1325 0.5325 ;
        RECT 4.0575 0.7125 4.1325 0.7875 ;
        RECT 3.0600 0.2025 3.1350 0.2775 ;
        RECT 2.1900 0.6525 2.2650 0.7275 ;
        RECT 2.1525 0.3300 2.2275 0.4050 ;
        RECT 1.3875 0.3150 1.4625 0.3900 ;
        RECT 1.3875 0.6525 1.4625 0.7275 ;
        LAYER M2 ;
        RECT 5.1825 0.4200 5.3025 0.5700 ;
        RECT 5.1075 0.4200 5.1825 0.9375 ;
        RECT 4.3500 0.8625 5.1075 0.9375 ;
        RECT 4.2750 0.2100 4.3500 0.9375 ;
        RECT 4.0425 0.2100 4.2750 0.2850 ;
        RECT 4.0125 0.7125 4.2750 0.7875 ;
        RECT 4.0425 0.4125 4.1475 0.5775 ;
        RECT 3.9675 0.1125 4.0425 0.2850 ;
        RECT 3.5025 0.4125 4.0425 0.4875 ;
        RECT 3.1350 0.1125 3.9675 0.1875 ;
        RECT 3.4275 0.4125 3.5025 0.7275 ;
        RECT 2.0700 0.6525 3.4275 0.7275 ;
        RECT 3.0600 0.1125 3.1350 0.3525 ;
        RECT 2.0700 0.3150 2.2650 0.4200 ;
        RECT 1.9950 0.3150 2.0700 0.7275 ;
        RECT 1.5075 0.6525 1.9950 0.7275 ;
        RECT 1.4325 0.3150 1.5075 0.7275 ;
        RECT 1.3425 0.3150 1.4325 0.3900 ;
        RECT 1.3425 0.6525 1.4325 0.7275 ;
    END
END FA1_0111


MACRO FA1_1000
    CLASS CORE ;
    FOREIGN FA1_1000 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.5700 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 3.4575 0.1500 3.5325 0.9000 ;
        RECT 3.4050 0.1500 3.4575 0.2325 ;
        RECT 3.4125 0.6675 3.4575 0.9000 ;
        END
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 3.0375 0.2700 3.0675 0.4200 ;
        RECT 2.9625 0.2700 3.0375 0.9375 ;
        RECT 2.4900 0.8625 2.9625 0.9375 ;
        VIA 3.0150 0.3450 VIA12_square ;
        VIA 3.0000 0.7950 VIA12_square ;
        END
    END CO
    PIN CI
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.9425 0.3750 2.0475 0.5925 ;
        RECT 1.5150 0.5175 1.9425 0.5925 ;
        RECT 1.4400 0.2625 1.5150 0.5925 ;
        RECT 1.2300 0.2625 1.4400 0.3375 ;
        RECT 1.0800 0.2625 1.2300 0.4350 ;
        RECT 0.8250 0.2625 1.0800 0.3375 ;
        VIA 1.9950 0.4575 VIA12_square ;
        VIA 1.1550 0.3825 VIA12_square ;
        END
    END CI
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.6650 0.3600 1.7625 0.4350 ;
        RECT 1.5900 0.1125 1.6650 0.4350 ;
        RECT 0.5850 0.1125 1.5900 0.1875 ;
        RECT 0.5100 0.1125 0.5850 0.4875 ;
        RECT 0.3600 0.4125 0.5100 0.4875 ;
        VIA 1.6800 0.3975 VIA12_square ;
        VIA 0.4725 0.4500 VIA12_square ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 2.3700 0.4725 2.5425 0.5775 ;
        RECT 2.2950 0.4725 2.3700 0.8925 ;
        RECT 1.5450 0.8175 2.2950 0.8925 ;
        RECT 1.4700 0.8175 1.5450 0.9375 ;
        RECT 0.9300 0.8625 1.4700 0.9375 ;
        RECT 0.8550 0.8175 0.9300 0.9375 ;
        RECT 0.7050 0.8175 0.8550 0.8925 ;
        VIA 2.4600 0.5250 VIA12_square ;
        VIA 1.5825 0.8550 VIA12_square ;
        VIA 0.8175 0.8550 VIA12_square ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 3.3000 -0.0750 3.5700 0.0750 ;
        RECT 3.1950 -0.0750 3.3000 0.2325 ;
        RECT 2.4750 -0.0750 3.1950 0.0750 ;
        RECT 2.3550 -0.0750 2.4750 0.1800 ;
        RECT 2.0325 -0.0750 2.3550 0.0750 ;
        RECT 1.9575 -0.0750 2.0325 0.2625 ;
        RECT 0.5850 -0.0750 1.9575 0.0750 ;
        RECT 0.4650 -0.0750 0.5850 0.1800 ;
        RECT 0.1425 -0.0750 0.4650 0.0750 ;
        RECT 0.0675 -0.0750 0.1425 0.3075 ;
        RECT 0.0000 -0.0750 0.0675 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 3.3075 0.9750 3.5700 1.1250 ;
        RECT 3.2025 0.7950 3.3075 1.1250 ;
        RECT 2.4750 0.9750 3.2025 1.1250 ;
        RECT 2.3550 0.8700 2.4750 1.1250 ;
        RECT 2.0550 0.9750 2.3550 1.1250 ;
        RECT 1.9350 0.8025 2.0550 1.1250 ;
        RECT 0.5625 0.9750 1.9350 1.1250 ;
        RECT 0.4875 0.7800 0.5625 1.1250 ;
        RECT 0.1425 0.9750 0.4875 1.1250 ;
        RECT 0.0675 0.7875 0.1425 1.1250 ;
        RECT 0.0000 0.9750 0.0675 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 3.4350 0.1575 3.4950 0.2175 ;
        RECT 3.4350 0.8175 3.4950 0.8775 ;
        RECT 3.3225 0.4800 3.3825 0.5400 ;
        RECT 3.2250 0.1425 3.2850 0.2025 ;
        RECT 3.2250 0.8250 3.2850 0.8850 ;
        RECT 3.1125 0.5175 3.1725 0.5775 ;
        RECT 3.0150 0.1575 3.0750 0.2175 ;
        RECT 3.0150 0.8250 3.0750 0.8850 ;
        RECT 2.8050 0.1950 2.8650 0.2550 ;
        RECT 2.8050 0.7800 2.8650 0.8400 ;
        RECT 2.7000 0.5025 2.7600 0.5625 ;
        RECT 2.5950 0.2100 2.6550 0.2700 ;
        RECT 2.5950 0.7800 2.6550 0.8400 ;
        RECT 2.4900 0.5100 2.5500 0.5700 ;
        RECT 2.3850 0.1200 2.4450 0.1800 ;
        RECT 2.3850 0.8700 2.4450 0.9300 ;
        RECT 2.2800 0.5100 2.3400 0.5700 ;
        RECT 2.1750 0.1950 2.2350 0.2550 ;
        RECT 2.1750 0.7875 2.2350 0.8475 ;
        RECT 2.0625 0.4200 2.1225 0.4800 ;
        RECT 1.9650 0.1725 2.0250 0.2325 ;
        RECT 1.9650 0.8250 2.0250 0.8850 ;
        RECT 1.8675 0.4200 1.9275 0.4800 ;
        RECT 1.6500 0.5100 1.7100 0.5700 ;
        RECT 1.4400 0.5100 1.5000 0.5700 ;
        RECT 1.3350 0.1950 1.3950 0.2550 ;
        RECT 1.3350 0.7800 1.3950 0.8400 ;
        RECT 1.1250 0.1575 1.1850 0.2175 ;
        RECT 1.1250 0.6825 1.1850 0.7425 ;
        RECT 1.0200 0.4725 1.0800 0.5325 ;
        RECT 0.9150 0.3000 0.9750 0.3600 ;
        RECT 0.9150 0.6450 0.9750 0.7050 ;
        RECT 0.8100 0.8400 0.8700 0.9000 ;
        RECT 0.6000 0.4275 0.6600 0.4875 ;
        RECT 0.4950 0.1200 0.5550 0.1800 ;
        RECT 0.4950 0.8325 0.5550 0.8925 ;
        RECT 0.3900 0.4275 0.4500 0.4875 ;
        RECT 0.2850 0.2550 0.3450 0.3150 ;
        RECT 0.2850 0.7200 0.3450 0.7800 ;
        RECT 0.1800 0.4800 0.2400 0.5400 ;
        RECT 0.0750 0.2025 0.1350 0.2625 ;
        RECT 0.0750 0.8325 0.1350 0.8925 ;
        LAYER M1 ;
        RECT 3.2700 0.3075 3.3825 0.5925 ;
        RECT 3.0675 0.4950 3.1950 0.6075 ;
        RECT 2.9625 0.6975 3.1275 0.9000 ;
        RECT 2.9625 0.1500 3.1125 0.4200 ;
        RECT 2.7375 0.4950 3.0675 0.5850 ;
        RECT 2.8125 0.1500 2.8875 0.3825 ;
        RECT 2.7375 0.6600 2.8875 0.9000 ;
        RECT 2.7300 0.1500 2.8125 0.3450 ;
        RECT 2.6325 0.4200 2.7375 0.5850 ;
        RECT 2.5725 0.7200 2.6625 0.8700 ;
        RECT 2.5800 0.1800 2.6550 0.3300 ;
        RECT 2.2575 0.2550 2.5800 0.3300 ;
        RECT 2.2575 0.7200 2.5725 0.7950 ;
        RECT 2.4225 0.4050 2.5575 0.6450 ;
        RECT 2.2725 0.4650 2.3475 0.6450 ;
        RECT 1.7175 0.5700 2.2725 0.6450 ;
        RECT 2.1525 0.1725 2.2575 0.3300 ;
        RECT 2.1525 0.7200 2.2575 0.8700 ;
        RECT 1.9425 0.4050 2.1675 0.4950 ;
        RECT 1.8225 0.4200 1.9425 0.4950 ;
        RECT 1.8075 0.1500 1.8825 0.3150 ;
        RECT 1.4025 0.1500 1.8075 0.2250 ;
        RECT 1.6425 0.3000 1.7175 0.6450 ;
        RECT 1.5525 0.7875 1.6650 0.9000 ;
        RECT 1.6125 0.3000 1.6425 0.3750 ;
        RECT 1.4775 0.4650 1.5525 0.9000 ;
        RECT 1.4400 0.4650 1.4775 0.6075 ;
        RECT 1.3650 0.1500 1.4025 0.3750 ;
        RECT 1.3650 0.6825 1.4025 0.8700 ;
        RECT 1.3275 0.1500 1.3650 0.8700 ;
        RECT 1.2900 0.3000 1.3275 0.7575 ;
        RECT 0.7350 0.1500 1.2150 0.2250 ;
        RECT 1.1100 0.3000 1.2150 0.5325 ;
        RECT 1.0500 0.6075 1.2150 0.8325 ;
        RECT 0.9900 0.4575 1.1100 0.5325 ;
        RECT 0.8850 0.3000 1.0050 0.3750 ;
        RECT 0.8850 0.6150 0.9750 0.7350 ;
        RECT 0.7350 0.8175 0.9000 0.9000 ;
        RECT 0.8100 0.3000 0.8850 0.7350 ;
        RECT 0.6600 0.1500 0.7350 0.3300 ;
        RECT 0.6600 0.5625 0.7350 0.9000 ;
        RECT 0.3450 0.4050 0.7050 0.4875 ;
        RECT 0.2550 0.2550 0.6600 0.3300 ;
        RECT 0.2400 0.5625 0.6600 0.6375 ;
        RECT 0.2175 0.7125 0.4125 0.8775 ;
        RECT 0.1650 0.4350 0.2400 0.6375 ;
        LAYER VIA1 ;
        RECT 3.2775 0.4125 3.3525 0.4875 ;
        RECT 2.7675 0.1650 2.8425 0.2400 ;
        RECT 2.7675 0.6975 2.8425 0.7725 ;
        RECT 2.6475 0.4575 2.7225 0.5325 ;
        RECT 1.8075 0.1950 1.8825 0.2700 ;
        RECT 1.0950 0.6750 1.1700 0.7500 ;
        RECT 0.8100 0.5100 0.8850 0.5850 ;
        RECT 0.2775 0.7125 0.3525 0.7875 ;
        LAYER M2 ;
        RECT 3.2175 0.4125 3.4275 0.4875 ;
        RECT 3.1425 0.1200 3.2175 0.4875 ;
        RECT 2.8875 0.1200 3.1425 0.1950 ;
        RECT 2.8125 0.1200 2.8875 0.7875 ;
        RECT 1.9275 0.1650 2.8125 0.2400 ;
        RECT 2.7300 0.6825 2.8125 0.7875 ;
        RECT 2.6325 0.3150 2.7375 0.5775 ;
        RECT 2.2050 0.3150 2.6325 0.3900 ;
        RECT 2.1300 0.3150 2.2050 0.7425 ;
        RECT 1.3650 0.6675 2.1300 0.7425 ;
        RECT 1.7625 0.1650 1.9275 0.2850 ;
        RECT 1.2900 0.5100 1.3650 0.7425 ;
        RECT 0.7350 0.5100 1.2900 0.5850 ;
        RECT 1.0500 0.6600 1.2150 0.7650 ;
        RECT 0.3675 0.6600 1.0500 0.7350 ;
        RECT 0.2625 0.6600 0.3675 0.8325 ;
    END
END FA1_1000


MACRO FA1_1001
    CLASS CORE ;
    FOREIGN FA1_1001 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.2500 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 5.1375 0.1500 5.2125 0.9000 ;
        RECT 5.1075 0.1500 5.1375 0.2775 ;
        RECT 5.0850 0.8250 5.1375 0.9000 ;
        END
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 4.6425 0.7275 4.7475 0.9375 ;
        RECT 4.2075 0.8625 4.6425 0.9375 ;
        VIA 4.6950 0.8175 VIA12_square ;
        END
    END CO
    PIN CI
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 2.0325 0.4950 2.7225 0.5700 ;
        RECT 1.9575 0.4125 2.0325 0.5700 ;
        RECT 1.6050 0.4125 1.9575 0.4875 ;
        RECT 1.4400 0.4125 1.6050 0.5475 ;
        VIA 2.6400 0.5325 VIA12_square ;
        VIA 1.5225 0.4950 VIA12_square ;
        END
    END CI
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 3.3975 0.3450 3.5100 0.6225 ;
        RECT 2.1825 0.3450 3.3975 0.4200 ;
        RECT 2.1075 0.2625 2.1825 0.4200 ;
        RECT 0.9975 0.2625 2.1075 0.3375 ;
        RECT 0.8925 0.2625 0.9975 0.5475 ;
        VIA 3.4500 0.5325 VIA12_square ;
        VIA 2.2200 0.3825 VIA12_square ;
        VIA 0.9450 0.4650 VIA12_square ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 3.7800 0.5100 3.9150 0.6150 ;
        RECT 3.7050 0.5100 3.7800 0.7875 ;
        RECT 2.0625 0.7125 3.7050 0.7875 ;
        RECT 1.9875 0.6450 2.0625 0.7875 ;
        RECT 1.2900 0.6450 1.9875 0.7200 ;
        RECT 1.1850 0.4575 1.2900 0.7875 ;
        RECT 0.4650 0.7125 1.1850 0.7875 ;
        RECT 0.3900 0.4125 0.4650 0.7875 ;
        RECT 0.2850 0.4125 0.3900 0.4875 ;
        VIA 3.8325 0.5625 VIA12_square ;
        VIA 2.1450 0.7500 VIA12_square ;
        VIA 1.2375 0.5400 VIA12_square ;
        VIA 0.3675 0.4500 VIA12_square ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 5.0025 -0.0750 5.2500 0.0750 ;
        RECT 4.8675 -0.0750 5.0025 0.1875 ;
        RECT 3.9450 -0.0750 4.8675 0.0750 ;
        RECT 3.8250 -0.0750 3.9450 0.1800 ;
        RECT 3.5250 -0.0750 3.8250 0.0750 ;
        RECT 3.4050 -0.0750 3.5250 0.1800 ;
        RECT 3.1050 -0.0750 3.4050 0.0750 ;
        RECT 2.9850 -0.0750 3.1050 0.1800 ;
        RECT 2.6700 -0.0750 2.9850 0.0750 ;
        RECT 2.5950 -0.0750 2.6700 0.2475 ;
        RECT 1.0050 -0.0750 2.5950 0.0750 ;
        RECT 0.8850 -0.0750 1.0050 0.1800 ;
        RECT 0.5850 -0.0750 0.8850 0.0750 ;
        RECT 0.4650 -0.0750 0.5850 0.1800 ;
        RECT 0.1575 -0.0750 0.4650 0.0750 ;
        RECT 0.0525 -0.0750 0.1575 0.3150 ;
        RECT 0.0000 -0.0750 0.0525 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 4.9725 0.9750 5.2500 1.1250 ;
        RECT 4.8975 0.8325 4.9725 1.1250 ;
        RECT 3.9450 0.9750 4.8975 1.1250 ;
        RECT 3.8250 0.8700 3.9450 1.1250 ;
        RECT 3.5250 0.9750 3.8250 1.1250 ;
        RECT 3.4050 0.8700 3.5250 1.1250 ;
        RECT 3.1050 0.9750 3.4050 1.1250 ;
        RECT 2.9850 0.8700 3.1050 1.1250 ;
        RECT 2.6850 0.9750 2.9850 1.1250 ;
        RECT 2.5650 0.8025 2.6850 1.1250 ;
        RECT 0.9975 0.9750 2.5650 1.1250 ;
        RECT 0.8925 0.8250 0.9975 1.1250 ;
        RECT 0.5775 0.9750 0.8925 1.1250 ;
        RECT 0.4725 0.8250 0.5775 1.1250 ;
        RECT 0.1425 0.9750 0.4725 1.1250 ;
        RECT 0.0675 0.8025 0.1425 1.1250 ;
        RECT 0.0000 0.9750 0.0675 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 5.1150 0.1800 5.1750 0.2400 ;
        RECT 5.1150 0.8325 5.1750 0.8925 ;
        RECT 5.0025 0.4800 5.0625 0.5400 ;
        RECT 4.9050 0.1275 4.9650 0.1875 ;
        RECT 4.9050 0.8625 4.9650 0.9225 ;
        RECT 4.8075 0.4950 4.8675 0.5550 ;
        RECT 4.6950 0.1800 4.7550 0.2400 ;
        RECT 4.6950 0.8325 4.7550 0.8925 ;
        RECT 4.4850 0.1575 4.5450 0.2175 ;
        RECT 4.4850 0.8175 4.5450 0.8775 ;
        RECT 4.3725 0.4800 4.4325 0.5400 ;
        RECT 4.2750 0.3000 4.3350 0.3600 ;
        RECT 4.2750 0.6675 4.3350 0.7275 ;
        RECT 4.1700 0.4800 4.2300 0.5400 ;
        RECT 4.0650 0.2100 4.1250 0.2700 ;
        RECT 4.0650 0.7500 4.1250 0.8100 ;
        RECT 3.9525 0.4800 4.0125 0.5400 ;
        RECT 3.8550 0.1200 3.9150 0.1800 ;
        RECT 3.8550 0.8700 3.9150 0.9300 ;
        RECT 3.7500 0.4800 3.8100 0.5400 ;
        RECT 3.6450 0.2550 3.7050 0.3150 ;
        RECT 3.6450 0.7350 3.7050 0.7950 ;
        RECT 3.5400 0.4800 3.6000 0.5400 ;
        RECT 3.4350 0.1200 3.4950 0.1800 ;
        RECT 3.4350 0.8700 3.4950 0.9300 ;
        RECT 3.3300 0.4800 3.3900 0.5400 ;
        RECT 3.2250 0.2250 3.2850 0.2850 ;
        RECT 3.2250 0.7350 3.2850 0.7950 ;
        RECT 3.1125 0.4950 3.1725 0.5550 ;
        RECT 3.0150 0.1200 3.0750 0.1800 ;
        RECT 3.0150 0.8700 3.0750 0.9300 ;
        RECT 2.9100 0.4950 2.9700 0.5550 ;
        RECT 2.8050 0.1650 2.8650 0.2250 ;
        RECT 2.8050 0.7500 2.8650 0.8100 ;
        RECT 2.5950 0.1575 2.6550 0.2175 ;
        RECT 2.5950 0.8325 2.6550 0.8925 ;
        RECT 2.4975 0.4950 2.5575 0.5550 ;
        RECT 2.2725 0.5100 2.3325 0.5700 ;
        RECT 2.0775 0.5550 2.1375 0.6150 ;
        RECT 1.9650 0.1650 2.0250 0.2250 ;
        RECT 1.9650 0.7950 2.0250 0.8550 ;
        RECT 1.7550 0.3000 1.8150 0.3600 ;
        RECT 1.7550 0.7350 1.8150 0.7950 ;
        RECT 1.6425 0.4800 1.7025 0.5400 ;
        RECT 1.5450 0.1575 1.6050 0.2175 ;
        RECT 1.5450 0.6825 1.6050 0.7425 ;
        RECT 1.4400 0.4800 1.5000 0.5400 ;
        RECT 1.3350 0.3000 1.3950 0.3600 ;
        RECT 1.3350 0.8325 1.3950 0.8925 ;
        RECT 1.2300 0.4950 1.2900 0.5550 ;
        RECT 1.0200 0.4725 1.0800 0.5325 ;
        RECT 0.9150 0.1200 0.9750 0.1800 ;
        RECT 0.9150 0.8475 0.9750 0.9075 ;
        RECT 0.8100 0.4725 0.8700 0.5325 ;
        RECT 0.7050 0.2550 0.7650 0.3150 ;
        RECT 0.7050 0.7575 0.7650 0.8175 ;
        RECT 0.6000 0.4725 0.6600 0.5325 ;
        RECT 0.4950 0.1200 0.5550 0.1800 ;
        RECT 0.4950 0.8475 0.5550 0.9075 ;
        RECT 0.3900 0.4800 0.4500 0.5400 ;
        RECT 0.2850 0.2550 0.3450 0.3150 ;
        RECT 0.2850 0.7575 0.3450 0.8175 ;
        RECT 0.1800 0.4800 0.2400 0.5400 ;
        RECT 0.0750 0.2325 0.1350 0.2925 ;
        RECT 0.0750 0.8325 0.1350 0.8925 ;
        LAYER M1 ;
        RECT 4.9875 0.3525 5.0625 0.7200 ;
        RECT 4.8300 0.3675 4.9125 0.7275 ;
        RECT 4.8225 0.4575 4.8300 0.7275 ;
        RECT 4.8075 0.4575 4.8225 0.6525 ;
        RECT 4.7550 0.1500 4.7850 0.2700 ;
        RECT 4.7325 0.8250 4.7850 0.9000 ;
        RECT 4.7325 0.1500 4.7550 0.3525 ;
        RECT 4.6800 0.1500 4.7325 0.9000 ;
        RECT 4.6575 0.2925 4.6800 0.9000 ;
        RECT 4.5075 0.3000 4.5825 0.7200 ;
        RECT 4.1250 0.1500 4.5750 0.2250 ;
        RECT 4.4625 0.7950 4.5675 0.9000 ;
        RECT 4.2450 0.3000 4.5075 0.3750 ;
        RECT 4.3575 0.6450 4.5075 0.7200 ;
        RECT 4.1325 0.8250 4.4625 0.9000 ;
        RECT 4.0875 0.4500 4.4325 0.5700 ;
        RECT 4.2525 0.6450 4.3575 0.7500 ;
        RECT 4.0575 0.7200 4.1325 0.9000 ;
        RECT 4.0500 0.1500 4.1250 0.3300 ;
        RECT 2.8725 0.7200 4.0575 0.7950 ;
        RECT 3.3075 0.2550 4.0500 0.3300 ;
        RECT 3.7500 0.4500 4.0125 0.6150 ;
        RECT 3.3300 0.4500 3.6000 0.5850 ;
        RECT 3.2025 0.2025 3.3075 0.3300 ;
        RECT 2.8950 0.2550 3.2025 0.3300 ;
        RECT 2.6925 0.4800 3.2025 0.5700 ;
        RECT 2.7750 0.1500 2.8950 0.3300 ;
        RECT 2.7975 0.7200 2.8725 0.8400 ;
        RECT 2.4375 0.4650 2.6925 0.5700 ;
        RECT 2.3250 0.1500 2.4900 0.2325 ;
        RECT 2.2575 0.3450 2.3625 0.6450 ;
        RECT 2.0025 0.1500 2.3250 0.2250 ;
        RECT 2.1825 0.8025 2.2725 0.9000 ;
        RECT 2.1375 0.3450 2.2575 0.4200 ;
        RECT 2.1075 0.5250 2.1825 0.9000 ;
        RECT 2.0775 0.5250 2.1075 0.6450 ;
        RECT 2.0025 0.7650 2.0325 0.8850 ;
        RECT 1.9275 0.1500 2.0025 0.8850 ;
        RECT 1.7775 0.3000 1.8525 0.9000 ;
        RECT 1.3050 0.3000 1.7775 0.3750 ;
        RECT 1.7475 0.6975 1.7775 0.9000 ;
        RECT 1.6500 0.8175 1.7475 0.9000 ;
        RECT 1.4400 0.4500 1.7025 0.5850 ;
        RECT 1.3050 0.8250 1.6500 0.9000 ;
        RECT 1.1550 0.1500 1.6350 0.2250 ;
        RECT 1.5150 0.6675 1.6350 0.7425 ;
        RECT 1.4400 0.6675 1.5150 0.7500 ;
        RECT 0.7875 0.6750 1.4400 0.7500 ;
        RECT 1.1550 0.4500 1.3650 0.6000 ;
        RECT 1.0800 0.1500 1.1550 0.3375 ;
        RECT 0.7875 0.2625 1.0800 0.3375 ;
        RECT 0.5550 0.4275 1.0800 0.5700 ;
        RECT 0.6825 0.2100 0.7875 0.3375 ;
        RECT 0.6825 0.6750 0.7875 0.8400 ;
        RECT 0.3675 0.2625 0.6825 0.3375 ;
        RECT 0.3675 0.6750 0.6825 0.7500 ;
        RECT 0.1575 0.4125 0.4500 0.5850 ;
        RECT 0.2625 0.2100 0.3675 0.3375 ;
        RECT 0.2625 0.6750 0.3675 0.8400 ;
        LAYER VIA1 ;
        RECT 4.9875 0.4125 5.0625 0.4875 ;
        RECT 4.8225 0.6075 4.8975 0.6825 ;
        RECT 4.5075 0.4125 4.5825 0.4875 ;
        RECT 4.1325 0.4725 4.2075 0.5475 ;
        RECT 2.3700 0.1575 2.4450 0.2325 ;
        RECT 1.7325 0.8175 1.8075 0.8925 ;
        LAYER M2 ;
        RECT 4.3575 0.4125 5.1075 0.4875 ;
        RECT 4.8225 0.5625 4.8975 0.8100 ;
        RECT 4.2075 0.5625 4.8225 0.6375 ;
        RECT 4.2825 0.1425 4.3575 0.4875 ;
        RECT 2.4900 0.1425 4.2825 0.2175 ;
        RECT 4.1325 0.3975 4.2075 0.7875 ;
        RECT 4.0200 0.7125 4.1325 0.7875 ;
        RECT 3.9450 0.7125 4.0200 0.9375 ;
        RECT 1.8525 0.8625 3.9450 0.9375 ;
        RECT 2.3250 0.1425 2.4900 0.2475 ;
        RECT 1.6875 0.8025 1.8525 0.9375 ;
    END
END FA1_1001


MACRO FA1_1010
    CLASS CORE ;
    FOREIGN FA1_1010 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.5700 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 3.4575 0.2175 3.5325 0.8325 ;
        RECT 3.4275 0.2175 3.4575 0.3825 ;
        RECT 3.4275 0.6675 3.4575 0.8325 ;
        END
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 3.0375 0.2700 3.0675 0.4200 ;
        RECT 2.9625 0.2700 3.0375 0.9375 ;
        RECT 2.4900 0.8625 2.9625 0.9375 ;
        VIA 3.0150 0.3450 VIA12_square ;
        VIA 3.0000 0.7950 VIA12_square ;
        END
    END CO
    PIN CI
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.9425 0.3750 2.0475 0.5925 ;
        RECT 1.5150 0.5175 1.9425 0.5925 ;
        RECT 1.4400 0.2625 1.5150 0.5925 ;
        RECT 1.2300 0.2625 1.4400 0.3375 ;
        RECT 1.0800 0.2625 1.2300 0.4350 ;
        RECT 0.8250 0.2625 1.0800 0.3375 ;
        VIA 1.9950 0.4575 VIA12_square ;
        VIA 1.1550 0.3825 VIA12_square ;
        END
    END CI
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.6650 0.3600 1.7625 0.4350 ;
        RECT 1.5900 0.1125 1.6650 0.4350 ;
        RECT 0.5850 0.1125 1.5900 0.1875 ;
        RECT 0.5100 0.1125 0.5850 0.4875 ;
        RECT 0.3600 0.4125 0.5100 0.4875 ;
        VIA 1.6800 0.3975 VIA12_square ;
        VIA 0.4725 0.4500 VIA12_square ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 2.3700 0.4725 2.5425 0.5775 ;
        RECT 2.2950 0.4725 2.3700 0.8925 ;
        RECT 1.5450 0.8175 2.2950 0.8925 ;
        RECT 1.4700 0.8175 1.5450 0.9375 ;
        RECT 0.9300 0.8625 1.4700 0.9375 ;
        RECT 0.8550 0.8175 0.9300 0.9375 ;
        RECT 0.7050 0.8175 0.8550 0.8925 ;
        VIA 2.4600 0.5250 VIA12_square ;
        VIA 1.5825 0.8550 VIA12_square ;
        VIA 0.8175 0.8550 VIA12_square ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 3.3225 -0.0750 3.5700 0.0750 ;
        RECT 3.1875 -0.0750 3.3225 0.2400 ;
        RECT 2.4750 -0.0750 3.1875 0.0750 ;
        RECT 2.3550 -0.0750 2.4750 0.1800 ;
        RECT 2.0325 -0.0750 2.3550 0.0750 ;
        RECT 1.9575 -0.0750 2.0325 0.2625 ;
        RECT 0.5850 -0.0750 1.9575 0.0750 ;
        RECT 0.4650 -0.0750 0.5850 0.1800 ;
        RECT 0.1425 -0.0750 0.4650 0.0750 ;
        RECT 0.0675 -0.0750 0.1425 0.3075 ;
        RECT 0.0000 -0.0750 0.0675 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 3.3075 0.9750 3.5700 1.1250 ;
        RECT 3.2025 0.7200 3.3075 1.1250 ;
        RECT 2.4750 0.9750 3.2025 1.1250 ;
        RECT 2.3550 0.8700 2.4750 1.1250 ;
        RECT 2.0550 0.9750 2.3550 1.1250 ;
        RECT 1.9350 0.8025 2.0550 1.1250 ;
        RECT 0.5625 0.9750 1.9350 1.1250 ;
        RECT 0.4875 0.7800 0.5625 1.1250 ;
        RECT 0.1425 0.9750 0.4875 1.1250 ;
        RECT 0.0675 0.7875 0.1425 1.1250 ;
        RECT 0.0000 0.9750 0.0675 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 3.4350 0.2700 3.4950 0.3300 ;
        RECT 3.4350 0.7200 3.4950 0.7800 ;
        RECT 3.3225 0.4950 3.3825 0.5550 ;
        RECT 3.2250 0.1800 3.2850 0.2400 ;
        RECT 3.2250 0.7500 3.2850 0.8100 ;
        RECT 3.1200 0.5175 3.1800 0.5775 ;
        RECT 3.0150 0.2325 3.0750 0.2925 ;
        RECT 3.0150 0.7575 3.0750 0.8175 ;
        RECT 2.8050 0.1950 2.8650 0.2550 ;
        RECT 2.8050 0.7800 2.8650 0.8400 ;
        RECT 2.7000 0.5025 2.7600 0.5625 ;
        RECT 2.5950 0.2100 2.6550 0.2700 ;
        RECT 2.5950 0.7800 2.6550 0.8400 ;
        RECT 2.4900 0.5100 2.5500 0.5700 ;
        RECT 2.3850 0.1200 2.4450 0.1800 ;
        RECT 2.3850 0.8700 2.4450 0.9300 ;
        RECT 2.2800 0.5100 2.3400 0.5700 ;
        RECT 2.1750 0.1950 2.2350 0.2550 ;
        RECT 2.1750 0.7875 2.2350 0.8475 ;
        RECT 2.0625 0.4200 2.1225 0.4800 ;
        RECT 1.9650 0.1725 2.0250 0.2325 ;
        RECT 1.9650 0.8250 2.0250 0.8850 ;
        RECT 1.8675 0.4200 1.9275 0.4800 ;
        RECT 1.6500 0.5100 1.7100 0.5700 ;
        RECT 1.4400 0.5100 1.5000 0.5700 ;
        RECT 1.3350 0.1950 1.3950 0.2550 ;
        RECT 1.3350 0.7800 1.3950 0.8400 ;
        RECT 1.1250 0.1575 1.1850 0.2175 ;
        RECT 1.1250 0.6825 1.1850 0.7425 ;
        RECT 1.0200 0.4725 1.0800 0.5325 ;
        RECT 0.9150 0.3000 0.9750 0.3600 ;
        RECT 0.9150 0.6450 0.9750 0.7050 ;
        RECT 0.8100 0.8400 0.8700 0.9000 ;
        RECT 0.6000 0.4275 0.6600 0.4875 ;
        RECT 0.4950 0.1200 0.5550 0.1800 ;
        RECT 0.4950 0.8325 0.5550 0.8925 ;
        RECT 0.3900 0.4275 0.4500 0.4875 ;
        RECT 0.2850 0.2550 0.3450 0.3150 ;
        RECT 0.2850 0.7200 0.3450 0.7800 ;
        RECT 0.1800 0.4800 0.2400 0.5400 ;
        RECT 0.0750 0.2025 0.1350 0.2625 ;
        RECT 0.0750 0.8325 0.1350 0.8925 ;
        LAYER M1 ;
        RECT 3.3525 0.4500 3.3825 0.6000 ;
        RECT 3.2775 0.3150 3.3525 0.6000 ;
        RECT 3.2175 0.3150 3.2775 0.4200 ;
        RECT 3.0675 0.4950 3.2025 0.6075 ;
        RECT 2.9625 0.6975 3.1275 0.9000 ;
        RECT 2.9625 0.1500 3.1125 0.4200 ;
        RECT 2.7375 0.4950 3.0675 0.5850 ;
        RECT 2.8125 0.1500 2.8875 0.3825 ;
        RECT 2.7375 0.6600 2.8875 0.9000 ;
        RECT 2.7300 0.1500 2.8125 0.3450 ;
        RECT 2.6325 0.4200 2.7375 0.5850 ;
        RECT 2.5725 0.7200 2.6625 0.8700 ;
        RECT 2.5800 0.1800 2.6550 0.3300 ;
        RECT 2.2575 0.2550 2.5800 0.3300 ;
        RECT 2.2575 0.7200 2.5725 0.7950 ;
        RECT 2.4225 0.4050 2.5575 0.6450 ;
        RECT 2.2725 0.4650 2.3475 0.6450 ;
        RECT 1.7175 0.5700 2.2725 0.6450 ;
        RECT 2.1525 0.1725 2.2575 0.3300 ;
        RECT 2.1525 0.7200 2.2575 0.8700 ;
        RECT 1.9425 0.4050 2.1675 0.4950 ;
        RECT 1.8225 0.4200 1.9425 0.4950 ;
        RECT 1.8075 0.1500 1.8825 0.3150 ;
        RECT 1.4025 0.1500 1.8075 0.2250 ;
        RECT 1.6425 0.3000 1.7175 0.6450 ;
        RECT 1.5525 0.7875 1.6650 0.9000 ;
        RECT 1.6125 0.3000 1.6425 0.3750 ;
        RECT 1.4775 0.4650 1.5525 0.9000 ;
        RECT 1.4400 0.4650 1.4775 0.6075 ;
        RECT 1.3650 0.1500 1.4025 0.3750 ;
        RECT 1.3650 0.6825 1.4025 0.8700 ;
        RECT 1.3275 0.1500 1.3650 0.8700 ;
        RECT 1.2900 0.3000 1.3275 0.7575 ;
        RECT 0.7350 0.1500 1.2150 0.2250 ;
        RECT 1.1100 0.3000 1.2150 0.5325 ;
        RECT 1.0500 0.6075 1.2150 0.8325 ;
        RECT 0.9900 0.4575 1.1100 0.5325 ;
        RECT 0.8850 0.3000 1.0050 0.3750 ;
        RECT 0.8850 0.6150 0.9750 0.7350 ;
        RECT 0.7350 0.8175 0.9000 0.9000 ;
        RECT 0.8100 0.3000 0.8850 0.7350 ;
        RECT 0.6600 0.1500 0.7350 0.3300 ;
        RECT 0.6600 0.5625 0.7350 0.9000 ;
        RECT 0.3450 0.4050 0.7050 0.4875 ;
        RECT 0.2550 0.2550 0.6600 0.3300 ;
        RECT 0.2400 0.5625 0.6600 0.6375 ;
        RECT 0.2175 0.7125 0.4125 0.8775 ;
        RECT 0.1650 0.4350 0.2400 0.6375 ;
        LAYER VIA1 ;
        RECT 3.2775 0.4125 3.3525 0.4875 ;
        RECT 2.7675 0.1650 2.8425 0.2400 ;
        RECT 2.7675 0.6975 2.8425 0.7725 ;
        RECT 2.6475 0.4575 2.7225 0.5325 ;
        RECT 1.8075 0.1950 1.8825 0.2700 ;
        RECT 1.0950 0.6750 1.1700 0.7500 ;
        RECT 0.8100 0.5100 0.8850 0.5850 ;
        RECT 0.2775 0.7125 0.3525 0.7875 ;
        LAYER M2 ;
        RECT 3.2175 0.4125 3.4275 0.4875 ;
        RECT 3.1425 0.1200 3.2175 0.4875 ;
        RECT 2.8875 0.1200 3.1425 0.1950 ;
        RECT 2.8125 0.1200 2.8875 0.7875 ;
        RECT 1.9275 0.1650 2.8125 0.2400 ;
        RECT 2.7300 0.6825 2.8125 0.7875 ;
        RECT 2.6325 0.3150 2.7375 0.5775 ;
        RECT 2.2050 0.3150 2.6325 0.3900 ;
        RECT 2.1300 0.3150 2.2050 0.7425 ;
        RECT 1.3650 0.6675 2.1300 0.7425 ;
        RECT 1.7625 0.1650 1.9275 0.2850 ;
        RECT 1.2900 0.5100 1.3650 0.7425 ;
        RECT 0.7350 0.5100 1.2900 0.5850 ;
        RECT 1.0500 0.6600 1.2150 0.7650 ;
        RECT 0.3675 0.6600 1.0500 0.7350 ;
        RECT 0.2625 0.6600 0.3675 0.8325 ;
    END
END FA1_1010


MACRO FILL16_0010
    CLASS CORE ;
    FOREIGN FILL16_0010 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.3600 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.0000 -0.0750 3.3600 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.0000 0.9750 3.3600 1.1250 ;
        END
    END VDD
END FILL16_0010


MACRO FILL2_0010
    CLASS CORE ;
    FOREIGN FILL2_0010 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.4200 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.0000 -0.0750 0.4200 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.0000 0.9750 0.4200 1.1250 ;
        END
    END VDD
END FILL2_0010


MACRO FILL32_0010
    CLASS CORE ;
    FOREIGN FILL32_0010 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.7200 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.0000 -0.0750 6.7200 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.0000 0.9750 6.7200 1.1250 ;
        END
    END VDD
END FILL32_0010


MACRO FILL3_0010
    CLASS CORE ;
    FOREIGN FILL3_0010 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.6300 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.0000 -0.0750 0.6300 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.0000 0.9750 0.6300 1.1250 ;
        END
    END VDD
END FILL3_0010


MACRO FILL4_0010
    CLASS CORE ;
    FOREIGN FILL4_0010 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.8400 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.0000 -0.0750 0.8400 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.0000 0.9750 0.8400 1.1250 ;
        END
    END VDD
END FILL4_0010


MACRO FILL64_0010
    CLASS CORE ;
    FOREIGN FILL64_0010 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.4400 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.0000 -0.0750 13.4400 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.0000 0.9750 13.4400 1.1250 ;
        END
    END VDD
END FILL64_0010


MACRO FILL8_0010
    CLASS CORE ;
    FOREIGN FILL8_0010 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.6800 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.0000 -0.0750 1.6800 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.0000 0.9750 1.6800 1.1250 ;
        END
    END VDD
END FILL8_0010


MACRO HA1_0011
    CLASS CORE ;
    FOREIGN HA1_0011 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.1500 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 3.0375 0.3075 3.1125 0.7425 ;
        RECT 2.8725 0.3075 3.0375 0.3825 ;
        RECT 2.8725 0.6675 3.0375 0.7425 ;
        RECT 2.7975 0.2175 2.8725 0.3825 ;
        RECT 2.7975 0.6675 2.8725 0.8325 ;
        END
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.2775 0.2175 0.3525 0.3900 ;
        RECT 0.2775 0.6675 0.3525 0.8325 ;
        RECT 0.1125 0.3150 0.2775 0.3900 ;
        RECT 0.1125 0.6675 0.2775 0.7425 ;
        RECT 0.0375 0.3150 0.1125 0.7425 ;
        END
    END CO
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 2.3775 0.3375 2.5725 0.4425 ;
        RECT 2.3025 0.3375 2.3775 0.5700 ;
        RECT 1.9425 0.4950 2.3025 0.5700 ;
        RECT 1.8600 0.4650 1.9425 0.5700 ;
        RECT 1.7775 0.4650 1.8600 0.6375 ;
        RECT 1.1925 0.5625 1.7775 0.6375 ;
        RECT 1.0275 0.5625 1.1925 0.6450 ;
        VIA 2.4975 0.3900 VIA12_square ;
        VIA 1.8600 0.5100 VIA12_square ;
        VIA 1.1100 0.6075 VIA12_square ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.7950 0.4125 1.2600 0.4875 ;
        VIA 0.9375 0.4500 VIA12_square ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 3.1050 -0.0750 3.1500 0.0750 ;
        RECT 2.9850 -0.0750 3.1050 0.2325 ;
        RECT 2.6850 -0.0750 2.9850 0.0750 ;
        RECT 2.5800 -0.0750 2.6850 0.2250 ;
        RECT 1.6350 -0.0750 2.5800 0.0750 ;
        RECT 1.5150 -0.0750 1.6350 0.1800 ;
        RECT 1.2000 -0.0750 1.5150 0.0750 ;
        RECT 1.1100 -0.0750 1.2000 0.3000 ;
        RECT 0.5850 -0.0750 1.1100 0.0750 ;
        RECT 0.4650 -0.0750 0.5850 0.1875 ;
        RECT 0.1575 -0.0750 0.4650 0.0750 ;
        RECT 0.0525 -0.0750 0.1575 0.2400 ;
        RECT 0.0000 -0.0750 0.0525 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 3.1050 0.9750 3.1500 1.1250 ;
        RECT 2.9850 0.8175 3.1050 1.1250 ;
        RECT 2.6775 0.9750 2.9850 1.1250 ;
        RECT 2.5725 0.6825 2.6775 1.1250 ;
        RECT 1.4250 0.9750 2.5725 1.1250 ;
        RECT 1.3050 0.8700 1.4250 1.1250 ;
        RECT 0.9825 0.9750 1.3050 1.1250 ;
        RECT 0.9075 0.7500 0.9825 1.1250 ;
        RECT 0.5850 0.9750 0.9075 1.1250 ;
        RECT 0.4650 0.8700 0.5850 1.1250 ;
        RECT 0.1650 0.9750 0.4650 1.1250 ;
        RECT 0.0450 0.8175 0.1650 1.1250 ;
        RECT 0.0000 0.9750 0.0450 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 3.0150 0.1575 3.0750 0.2175 ;
        RECT 3.0150 0.8325 3.0750 0.8925 ;
        RECT 2.9025 0.4875 2.9625 0.5475 ;
        RECT 2.8050 0.2700 2.8650 0.3300 ;
        RECT 2.8050 0.7200 2.8650 0.7800 ;
        RECT 2.7000 0.4875 2.7600 0.5475 ;
        RECT 2.5950 0.1350 2.6550 0.1950 ;
        RECT 2.5950 0.7050 2.6550 0.7650 ;
        RECT 2.5950 0.8700 2.6550 0.9300 ;
        RECT 2.4900 0.4650 2.5500 0.5250 ;
        RECT 2.3850 0.1575 2.4450 0.2175 ;
        RECT 2.3850 0.7275 2.4450 0.7875 ;
        RECT 2.1750 0.2250 2.2350 0.2850 ;
        RECT 2.1750 0.8250 2.2350 0.8850 ;
        RECT 2.0700 0.4875 2.1300 0.5475 ;
        RECT 1.9650 0.1725 2.0250 0.2325 ;
        RECT 1.9650 0.6600 2.0250 0.7200 ;
        RECT 1.8600 0.4650 1.9200 0.5250 ;
        RECT 1.7550 0.6600 1.8150 0.7200 ;
        RECT 1.6500 0.4125 1.7100 0.4725 ;
        RECT 1.5450 0.1200 1.6050 0.1800 ;
        RECT 1.5450 0.8250 1.6050 0.8850 ;
        RECT 1.4400 0.4125 1.5000 0.4725 ;
        RECT 1.4400 0.6525 1.5000 0.7125 ;
        RECT 1.3350 0.2400 1.3950 0.3000 ;
        RECT 1.3350 0.8700 1.3950 0.9300 ;
        RECT 1.2300 0.4350 1.2900 0.4950 ;
        RECT 1.1250 0.1950 1.1850 0.2550 ;
        RECT 1.1250 0.7875 1.1850 0.8475 ;
        RECT 1.0200 0.4350 1.0800 0.4950 ;
        RECT 0.9150 0.2625 0.9750 0.3225 ;
        RECT 0.9150 0.7875 0.9750 0.8475 ;
        RECT 0.8100 0.4350 0.8700 0.4950 ;
        RECT 0.7050 0.7275 0.7650 0.7875 ;
        RECT 0.6000 0.4950 0.6600 0.5550 ;
        RECT 0.4950 0.1200 0.5550 0.1800 ;
        RECT 0.4950 0.8700 0.5550 0.9300 ;
        RECT 0.3900 0.4800 0.4500 0.5400 ;
        RECT 0.2850 0.2700 0.3450 0.3300 ;
        RECT 0.2850 0.7200 0.3450 0.7800 ;
        RECT 0.1875 0.4950 0.2475 0.5550 ;
        RECT 0.0750 0.1575 0.1350 0.2175 ;
        RECT 0.0750 0.8325 0.1350 0.8925 ;
        LAYER M1 ;
        RECT 2.7375 0.4575 2.9625 0.5775 ;
        RECT 2.6325 0.4575 2.7375 0.6075 ;
        RECT 2.5500 0.3000 2.6550 0.3825 ;
        RECT 2.4600 0.3000 2.5500 0.5625 ;
        RECT 2.3850 0.1500 2.4750 0.2250 ;
        RECT 2.3850 0.6675 2.4600 0.8325 ;
        RECT 2.3775 0.1500 2.3850 0.8325 ;
        RECT 2.3100 0.1500 2.3775 0.7425 ;
        RECT 2.0400 0.4875 2.3100 0.5625 ;
        RECT 1.6200 0.8175 2.2650 0.9000 ;
        RECT 2.1300 0.1650 2.2350 0.4125 ;
        RECT 1.9200 0.6375 2.2200 0.7425 ;
        RECT 2.0400 0.3300 2.1300 0.4125 ;
        RECT 1.9425 0.1500 2.0550 0.2550 ;
        RECT 1.7850 0.1500 1.9425 0.2775 ;
        RECT 1.7850 0.3525 1.9350 0.5625 ;
        RECT 1.7250 0.6375 1.8375 0.7425 ;
        RECT 1.7100 0.6375 1.7250 0.7200 ;
        RECT 1.6350 0.2550 1.7100 0.7200 ;
        RECT 1.4175 0.2550 1.6350 0.3300 ;
        RECT 1.4175 0.6450 1.6350 0.7200 ;
        RECT 1.5150 0.7950 1.6200 0.9000 ;
        RECT 1.4175 0.4125 1.5300 0.5175 ;
        RECT 1.3125 0.2100 1.4175 0.3300 ;
        RECT 0.7800 0.4125 1.4175 0.4950 ;
        RECT 1.3425 0.6450 1.4175 0.7950 ;
        RECT 1.2000 0.7200 1.3425 0.7950 ;
        RECT 0.6750 0.5700 1.2375 0.6450 ;
        RECT 1.1175 0.7200 1.2000 0.8775 ;
        RECT 0.5250 0.2625 1.0050 0.3375 ;
        RECT 0.5250 0.7200 0.8025 0.7950 ;
        RECT 0.6000 0.4650 0.6750 0.6450 ;
        RECT 0.4500 0.2625 0.5250 0.7950 ;
        RECT 0.1875 0.4650 0.4500 0.5850 ;
        LAYER VIA1 ;
        RECT 2.6475 0.4950 2.7225 0.5700 ;
        RECT 2.1075 0.3300 2.1825 0.4050 ;
        RECT 2.1000 0.6450 2.1750 0.7200 ;
        RECT 1.8450 0.1650 1.9200 0.2400 ;
        RECT 1.6350 0.3150 1.7100 0.3900 ;
        LAYER M2 ;
        RECT 2.6475 0.1650 2.7225 0.6375 ;
        RECT 1.8000 0.1650 2.6475 0.2400 ;
        RECT 2.5275 0.5625 2.6475 0.6375 ;
        RECT 2.4525 0.5625 2.5275 0.7200 ;
        RECT 2.0550 0.6450 2.4525 0.7200 ;
        RECT 2.0550 0.3150 2.2275 0.4200 ;
        RECT 1.5750 0.3150 2.0550 0.3900 ;
    END
END HA1_0011


MACRO HA1_0111
    CLASS CORE ;
    FOREIGN HA1_0111 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.8300 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 4.1475 0.2625 4.4625 0.7425 ;
        VIA 4.3050 0.3225 VIA12_slot ;
        VIA 4.3050 0.6825 VIA12_slot ;
        END
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 0.3675 0.2625 0.6825 0.7275 ;
        VIA 0.5250 0.3225 VIA12_slot ;
        VIA 0.5250 0.6675 VIA12_slot ;
        END
    END CO
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 3.6975 0.4500 3.8475 0.5550 ;
        RECT 2.1975 0.4800 3.6975 0.5550 ;
        RECT 2.1225 0.4125 2.1975 0.5550 ;
        RECT 1.6575 0.4125 2.1225 0.4875 ;
        RECT 1.5375 0.3075 1.6575 0.4875 ;
        VIA 3.7725 0.5025 VIA12_square ;
        VIA 3.0450 0.5175 VIA12_square ;
        VIA 1.6050 0.3825 VIA12_square ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.4175 0.5625 1.8825 0.6375 ;
        RECT 1.3125 0.4650 1.4175 0.6375 ;
        VIA 1.3650 0.5475 VIA12_square ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 4.7625 -0.0750 4.8300 0.0750 ;
        RECT 4.6875 -0.0750 4.7625 0.3150 ;
        RECT 4.3650 -0.0750 4.6875 0.0750 ;
        RECT 4.2450 -0.0750 4.3650 0.1950 ;
        RECT 3.9450 -0.0750 4.2450 0.0750 ;
        RECT 3.8400 -0.0750 3.9450 0.2250 ;
        RECT 2.8650 -0.0750 3.8400 0.0750 ;
        RECT 2.7600 -0.0750 2.8650 0.2250 ;
        RECT 2.2650 -0.0750 2.7600 0.0750 ;
        RECT 2.1450 -0.0750 2.2650 0.1950 ;
        RECT 1.8225 -0.0750 2.1450 0.0750 ;
        RECT 1.7475 -0.0750 1.8225 0.2400 ;
        RECT 0.9975 -0.0750 1.7475 0.0750 ;
        RECT 0.8925 -0.0750 0.9975 0.2700 ;
        RECT 0.5850 -0.0750 0.8925 0.0750 ;
        RECT 0.4650 -0.0750 0.5850 0.1950 ;
        RECT 0.1425 -0.0750 0.4650 0.0750 ;
        RECT 0.0675 -0.0750 0.1425 0.3150 ;
        RECT 0.0000 -0.0750 0.0675 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 4.7775 0.9750 4.8300 1.1250 ;
        RECT 4.6725 0.6450 4.7775 1.1250 ;
        RECT 4.3575 0.9750 4.6725 1.1250 ;
        RECT 4.2525 0.8025 4.3575 1.1250 ;
        RECT 3.9450 0.9750 4.2525 1.1250 ;
        RECT 3.8250 0.6900 3.9450 1.1250 ;
        RECT 2.8950 0.9750 3.8250 1.1250 ;
        RECT 2.7750 0.8175 2.8950 1.1250 ;
        RECT 2.4675 0.9750 2.7750 1.1250 ;
        RECT 2.3625 0.7950 2.4675 1.1250 ;
        RECT 2.2650 0.9750 2.3625 1.1250 ;
        RECT 2.1450 0.7950 2.2650 1.1250 ;
        RECT 1.8300 0.9750 2.1450 1.1250 ;
        RECT 1.7400 0.7575 1.8300 1.1250 ;
        RECT 1.4250 0.9750 1.7400 1.1250 ;
        RECT 1.3050 0.8700 1.4250 1.1250 ;
        RECT 1.0050 0.9750 1.3050 1.1250 ;
        RECT 0.8850 0.8700 1.0050 1.1250 ;
        RECT 0.5775 0.9750 0.8850 1.1250 ;
        RECT 0.4725 0.8025 0.5775 1.1250 ;
        RECT 0.1425 0.9750 0.4725 1.1250 ;
        RECT 0.0675 0.6375 0.1425 1.1250 ;
        RECT 0.0000 0.9750 0.0675 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 4.6950 0.2250 4.7550 0.2850 ;
        RECT 4.6950 0.6675 4.7550 0.7275 ;
        RECT 4.6950 0.8325 4.7550 0.8925 ;
        RECT 4.5900 0.4800 4.6500 0.5400 ;
        RECT 4.4850 0.2250 4.5450 0.2850 ;
        RECT 4.4850 0.7575 4.5450 0.8175 ;
        RECT 4.3800 0.4800 4.4400 0.5400 ;
        RECT 4.2750 0.1275 4.3350 0.1875 ;
        RECT 4.2750 0.8325 4.3350 0.8925 ;
        RECT 4.1700 0.4800 4.2300 0.5400 ;
        RECT 4.0650 0.2250 4.1250 0.2850 ;
        RECT 4.0650 0.7575 4.1250 0.8175 ;
        RECT 3.9600 0.4800 4.0200 0.5400 ;
        RECT 3.8550 0.1350 3.9150 0.1950 ;
        RECT 3.8550 0.7050 3.9150 0.7650 ;
        RECT 3.8550 0.8700 3.9150 0.9300 ;
        RECT 3.7500 0.4650 3.8100 0.5250 ;
        RECT 3.6450 0.1575 3.7050 0.2175 ;
        RECT 3.6450 0.7425 3.7050 0.8025 ;
        RECT 3.4350 0.2550 3.4950 0.3150 ;
        RECT 3.4350 0.6525 3.4950 0.7125 ;
        RECT 3.3375 0.4725 3.3975 0.5325 ;
        RECT 3.2250 0.1650 3.2850 0.2250 ;
        RECT 3.2250 0.8250 3.2850 0.8850 ;
        RECT 3.1125 0.4950 3.1725 0.5550 ;
        RECT 3.0150 0.3075 3.0750 0.3675 ;
        RECT 3.0150 0.8100 3.0750 0.8700 ;
        RECT 2.9100 0.6450 2.9700 0.7050 ;
        RECT 2.8050 0.1350 2.8650 0.1950 ;
        RECT 2.8050 0.8325 2.8650 0.8925 ;
        RECT 2.7000 0.4725 2.7600 0.5325 ;
        RECT 2.5950 0.2325 2.6550 0.2925 ;
        RECT 2.5950 0.7950 2.6550 0.8550 ;
        RECT 2.4900 0.4725 2.5500 0.5325 ;
        RECT 2.3850 0.2775 2.4450 0.3375 ;
        RECT 2.3850 0.8250 2.4450 0.8850 ;
        RECT 2.2800 0.4575 2.3400 0.5175 ;
        RECT 2.1750 0.1275 2.2350 0.1875 ;
        RECT 2.1750 0.8175 2.2350 0.8775 ;
        RECT 2.0700 0.4575 2.1300 0.5175 ;
        RECT 1.9650 0.2775 2.0250 0.3375 ;
        RECT 1.9650 0.7350 2.0250 0.7950 ;
        RECT 1.8600 0.4575 1.9200 0.5175 ;
        RECT 1.7550 0.1500 1.8150 0.2100 ;
        RECT 1.7550 0.7950 1.8150 0.8550 ;
        RECT 1.6500 0.4125 1.7100 0.4725 ;
        RECT 1.5450 0.7275 1.6050 0.7875 ;
        RECT 1.4400 0.4950 1.5000 0.5550 ;
        RECT 1.3350 0.1875 1.3950 0.2475 ;
        RECT 1.3350 0.8700 1.3950 0.9300 ;
        RECT 1.2300 0.4950 1.2900 0.5550 ;
        RECT 1.1250 0.7275 1.1850 0.7875 ;
        RECT 1.0200 0.4800 1.0800 0.5400 ;
        RECT 0.9150 0.1800 0.9750 0.2400 ;
        RECT 0.9150 0.8700 0.9750 0.9300 ;
        RECT 0.8100 0.4650 0.8700 0.5250 ;
        RECT 0.7050 0.2250 0.7650 0.2850 ;
        RECT 0.7050 0.7575 0.7650 0.8175 ;
        RECT 0.6000 0.4650 0.6600 0.5250 ;
        RECT 0.4950 0.1275 0.5550 0.1875 ;
        RECT 0.4950 0.8325 0.5550 0.8925 ;
        RECT 0.3900 0.4650 0.4500 0.5250 ;
        RECT 0.2850 0.2250 0.3450 0.2850 ;
        RECT 0.2850 0.7575 0.3450 0.8175 ;
        RECT 0.1800 0.4650 0.2400 0.5250 ;
        RECT 0.0750 0.2250 0.1350 0.2850 ;
        RECT 0.0750 0.6675 0.1350 0.7275 ;
        RECT 0.0750 0.8325 0.1350 0.8925 ;
        LAYER M1 ;
        RECT 3.8850 0.4575 4.6800 0.5625 ;
        RECT 4.4625 0.1950 4.5675 0.3675 ;
        RECT 4.4775 0.6375 4.5525 0.8700 ;
        RECT 4.1325 0.6375 4.4775 0.7275 ;
        RECT 4.1475 0.2775 4.4625 0.3675 ;
        RECT 4.0425 0.1950 4.1475 0.3675 ;
        RECT 4.0575 0.6375 4.1325 0.8700 ;
        RECT 3.8100 0.3000 3.9375 0.3825 ;
        RECT 3.7350 0.3000 3.8100 0.5850 ;
        RECT 3.6600 0.1500 3.7350 0.2250 ;
        RECT 3.6600 0.6900 3.7200 0.8625 ;
        RECT 3.6375 0.1500 3.6600 0.8625 ;
        RECT 3.5850 0.1500 3.6375 0.7650 ;
        RECT 3.3075 0.4725 3.5850 0.5475 ;
        RECT 3.2925 0.8175 3.5250 0.9000 ;
        RECT 3.4350 0.1800 3.5100 0.3975 ;
        RECT 3.3525 0.6225 3.5025 0.7425 ;
        RECT 3.2100 0.3225 3.4350 0.3975 ;
        RECT 3.3000 0.6225 3.3525 0.7200 ;
        RECT 3.1650 0.1500 3.3300 0.2475 ;
        RECT 3.1875 0.6450 3.3000 0.7200 ;
        RECT 3.1575 0.7950 3.2925 0.9000 ;
        RECT 3.0975 0.4725 3.2025 0.5700 ;
        RECT 2.9700 0.1500 3.1650 0.2250 ;
        RECT 2.6625 0.3000 3.1050 0.3750 ;
        RECT 2.9100 0.4500 3.0975 0.5700 ;
        RECT 2.9775 0.6450 3.0825 0.9000 ;
        RECT 2.8350 0.6450 2.9775 0.7200 ;
        RECT 2.7600 0.4650 2.8350 0.7200 ;
        RECT 2.4975 0.4650 2.7600 0.5400 ;
        RECT 2.5725 0.6150 2.6850 0.9000 ;
        RECT 2.5875 0.1950 2.6625 0.3750 ;
        RECT 2.4225 0.2700 2.4975 0.7050 ;
        RECT 1.9350 0.2700 2.4225 0.3450 ;
        RECT 2.0325 0.6300 2.4225 0.7050 ;
        RECT 1.8825 0.4275 2.3475 0.5475 ;
        RECT 1.9575 0.6300 2.0325 0.8325 ;
        RECT 1.8075 0.4275 1.8825 0.6450 ;
        RECT 1.5375 0.5700 1.8075 0.6450 ;
        RECT 1.6275 0.3450 1.7325 0.4950 ;
        RECT 0.9300 0.7200 1.6350 0.7950 ;
        RECT 1.1025 0.3450 1.6275 0.4200 ;
        RECT 1.4700 0.4950 1.5375 0.6450 ;
        RECT 1.2000 0.4950 1.4700 0.6075 ;
        RECT 1.0725 0.1650 1.4250 0.2700 ;
        RECT 1.0125 0.3450 1.1025 0.5925 ;
        RECT 0.8550 0.4425 0.9300 0.7950 ;
        RECT 0.1500 0.4425 0.8550 0.5475 ;
        RECT 0.6825 0.1950 0.7875 0.3675 ;
        RECT 0.6975 0.6225 0.7725 0.8700 ;
        RECT 0.3525 0.6225 0.6975 0.7125 ;
        RECT 0.3675 0.2775 0.6825 0.3675 ;
        RECT 0.2625 0.1950 0.3675 0.3675 ;
        RECT 0.2775 0.6225 0.3525 0.8700 ;
        LAYER VIA1 ;
        RECT 3.9375 0.4725 4.0125 0.5475 ;
        RECT 3.3900 0.8175 3.4650 0.8925 ;
        RECT 3.3600 0.3225 3.4350 0.3975 ;
        RECT 3.2325 0.6450 3.3075 0.7200 ;
        RECT 3.2100 0.1575 3.2850 0.2325 ;
        RECT 2.5950 0.6600 2.6700 0.7350 ;
        RECT 2.4225 0.3225 2.4975 0.3975 ;
        RECT 1.1325 0.7200 1.2075 0.7950 ;
        RECT 1.1175 0.1800 1.1925 0.2550 ;
        LAYER M2 ;
        RECT 3.9975 0.4350 4.0275 0.5850 ;
        RECT 3.9225 0.2625 3.9975 0.7875 ;
        RECT 3.7350 0.2625 3.9225 0.3375 ;
        RECT 3.6075 0.7125 3.9225 0.7875 ;
        RECT 3.6600 0.1575 3.7350 0.3375 ;
        RECT 3.1350 0.1575 3.6600 0.2325 ;
        RECT 3.5325 0.7125 3.6075 0.9000 ;
        RECT 3.3150 0.8175 3.5325 0.9000 ;
        RECT 2.3475 0.3225 3.5100 0.3975 ;
        RECT 2.7075 0.6450 3.3825 0.7200 ;
        RECT 2.5575 0.6450 2.7075 0.7500 ;
        RECT 1.1925 0.1650 1.2375 0.2700 ;
        RECT 1.1925 0.6825 1.2225 0.8325 ;
        RECT 1.1175 0.1650 1.1925 0.8325 ;
        RECT 1.0725 0.1650 1.1175 0.2700 ;
    END
END HA1_0111


MACRO HA1_1000
    CLASS CORE ;
    FOREIGN HA1_1000 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.7300 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 2.6175 0.1500 2.6925 0.9000 ;
        RECT 2.5650 0.1500 2.6175 0.3825 ;
        RECT 2.5725 0.7950 2.6175 0.9000 ;
        END
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1125 0.6675 0.1575 0.9000 ;
        RECT 0.1125 0.2025 0.1425 0.3225 ;
        RECT 0.0375 0.2025 0.1125 0.9000 ;
        END
    END CO
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 2.2575 0.4050 2.3625 0.5550 ;
        RECT 1.6200 0.4800 2.2575 0.5550 ;
        RECT 1.5450 0.4800 1.6200 0.6375 ;
        RECT 0.8625 0.5625 1.5450 0.6375 ;
        VIA 2.3100 0.4800 VIA12_square ;
        VIA 1.6425 0.5175 VIA12_square ;
        VIA 0.9450 0.6000 VIA12_square ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.8550 0.4125 1.3200 0.4875 ;
        VIA 1.0950 0.4500 VIA12_square ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 2.4750 -0.0750 2.7300 0.0750 ;
        RECT 2.3700 -0.0750 2.4750 0.2250 ;
        RECT 1.4250 -0.0750 2.3700 0.0750 ;
        RECT 1.3050 -0.0750 1.4250 0.1800 ;
        RECT 0.9900 -0.0750 1.3050 0.0750 ;
        RECT 0.9000 -0.0750 0.9900 0.3000 ;
        RECT 0.3750 -0.0750 0.9000 0.0750 ;
        RECT 0.2550 -0.0750 0.3750 0.1875 ;
        RECT 0.0000 -0.0750 0.2550 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 2.4750 0.9750 2.7300 1.1250 ;
        RECT 2.3550 0.8700 2.4750 1.1250 ;
        RECT 1.2150 0.9750 2.3550 1.1250 ;
        RECT 1.0950 0.8700 1.2150 1.1250 ;
        RECT 0.7725 0.9750 1.0950 1.1250 ;
        RECT 0.6975 0.7800 0.7725 1.1250 ;
        RECT 0.3750 0.9750 0.6975 1.1250 ;
        RECT 0.2550 0.8700 0.3750 1.1250 ;
        RECT 0.0000 0.9750 0.2550 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 2.5950 0.1575 2.6550 0.2175 ;
        RECT 2.5950 0.8175 2.6550 0.8775 ;
        RECT 2.4825 0.5100 2.5425 0.5700 ;
        RECT 2.3850 0.1350 2.4450 0.1950 ;
        RECT 2.3850 0.8700 2.4450 0.9300 ;
        RECT 2.2725 0.4650 2.3325 0.5250 ;
        RECT 2.1750 0.1575 2.2350 0.2175 ;
        RECT 2.1750 0.8100 2.2350 0.8700 ;
        RECT 1.9650 0.2250 2.0250 0.2850 ;
        RECT 1.9650 0.8175 2.0250 0.8775 ;
        RECT 1.8600 0.4800 1.9200 0.5400 ;
        RECT 1.7550 0.1725 1.8150 0.2325 ;
        RECT 1.7550 0.6900 1.8150 0.7500 ;
        RECT 1.6500 0.4425 1.7100 0.5025 ;
        RECT 1.5450 0.6900 1.6050 0.7500 ;
        RECT 1.4325 0.4125 1.4925 0.4725 ;
        RECT 1.3350 0.1200 1.3950 0.1800 ;
        RECT 1.3350 0.8250 1.3950 0.8850 ;
        RECT 1.2300 0.4125 1.2900 0.4725 ;
        RECT 1.2300 0.6525 1.2900 0.7125 ;
        RECT 1.1250 0.2400 1.1850 0.3000 ;
        RECT 1.1250 0.8700 1.1850 0.9300 ;
        RECT 1.0200 0.4275 1.0800 0.4875 ;
        RECT 0.9150 0.1950 0.9750 0.2550 ;
        RECT 0.9150 0.8100 0.9750 0.8700 ;
        RECT 0.8100 0.4275 0.8700 0.4875 ;
        RECT 0.7050 0.2100 0.7650 0.2700 ;
        RECT 0.7050 0.8175 0.7650 0.8775 ;
        RECT 0.6075 0.4275 0.6675 0.4875 ;
        RECT 0.4950 0.8175 0.5550 0.8775 ;
        RECT 0.3900 0.4950 0.4500 0.5550 ;
        RECT 0.2850 0.1200 0.3450 0.1800 ;
        RECT 0.2850 0.8700 0.3450 0.9300 ;
        RECT 0.1875 0.4800 0.2475 0.5400 ;
        RECT 0.0750 0.2325 0.1350 0.2925 ;
        RECT 0.0750 0.8175 0.1350 0.8775 ;
        LAYER M1 ;
        RECT 2.4975 0.4800 2.5425 0.6000 ;
        RECT 2.4225 0.4800 2.4975 0.7950 ;
        RECT 2.3475 0.3000 2.4675 0.4050 ;
        RECT 2.3325 0.6900 2.4225 0.7950 ;
        RECT 2.2725 0.3000 2.3475 0.5700 ;
        RECT 2.1975 0.1500 2.2650 0.2250 ;
        RECT 2.1975 0.6750 2.2575 0.9000 ;
        RECT 2.1525 0.1500 2.1975 0.9000 ;
        RECT 2.1225 0.1500 2.1525 0.7425 ;
        RECT 1.8300 0.4800 2.1225 0.5550 ;
        RECT 1.9500 0.1800 2.0475 0.4050 ;
        RECT 1.9425 0.7950 2.0475 0.9000 ;
        RECT 1.8825 0.6300 2.0175 0.7200 ;
        RECT 1.8150 0.3300 1.9500 0.4050 ;
        RECT 1.4100 0.8250 1.9425 0.9000 ;
        RECT 1.8000 0.6300 1.8825 0.7500 ;
        RECT 1.5750 0.1500 1.8750 0.2550 ;
        RECT 1.7100 0.6450 1.8000 0.7500 ;
        RECT 1.7100 0.4650 1.7175 0.5700 ;
        RECT 1.5675 0.3300 1.7100 0.5700 ;
        RECT 1.5150 0.6450 1.6350 0.7500 ;
        RECT 1.4925 0.6450 1.5150 0.7200 ;
        RECT 1.4175 0.2550 1.4925 0.7200 ;
        RECT 1.2075 0.2550 1.4175 0.3375 ;
        RECT 1.2075 0.6450 1.4175 0.7200 ;
        RECT 1.3050 0.7950 1.4100 0.9000 ;
        RECT 1.2075 0.4125 1.3200 0.5175 ;
        RECT 1.1025 0.2100 1.2075 0.3375 ;
        RECT 0.5700 0.4125 1.2075 0.4875 ;
        RECT 1.1325 0.6450 1.2075 0.7950 ;
        RECT 0.9975 0.7200 1.1325 0.7950 ;
        RECT 0.4650 0.5625 1.0275 0.6375 ;
        RECT 0.8925 0.7200 0.9975 0.9000 ;
        RECT 0.6750 0.2025 0.7950 0.3375 ;
        RECT 0.3150 0.2625 0.6750 0.3375 ;
        RECT 0.4725 0.7200 0.5775 0.9000 ;
        RECT 0.3150 0.7200 0.4725 0.7950 ;
        RECT 0.3900 0.4650 0.4650 0.6375 ;
        RECT 0.2400 0.2625 0.3150 0.7950 ;
        RECT 0.1875 0.4500 0.2400 0.5700 ;
        LAYER VIA1 ;
        RECT 2.3775 0.7125 2.4525 0.7875 ;
        RECT 1.8975 0.3300 1.9725 0.4050 ;
        RECT 1.7700 0.6600 1.8450 0.7350 ;
        RECT 1.6800 0.1575 1.7550 0.2325 ;
        RECT 1.3725 0.2625 1.4475 0.3375 ;
        LAYER M2 ;
        RECT 1.8825 0.7125 2.5275 0.7875 ;
        RECT 1.5600 0.3300 2.0175 0.4050 ;
        RECT 1.7325 0.6450 1.8825 0.7875 ;
        RECT 1.6350 0.1125 1.8000 0.2475 ;
        RECT 0.7050 0.7125 1.7325 0.7875 ;
        RECT 0.7050 0.1125 1.6350 0.1875 ;
        RECT 1.4775 0.2625 1.5600 0.4050 ;
        RECT 1.3275 0.2625 1.4775 0.3375 ;
        RECT 0.6300 0.1125 0.7050 0.7875 ;
    END
END HA1_1000


MACRO HA1_1010
    CLASS CORE ;
    FOREIGN HA1_1010 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.7300 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 2.6175 0.2175 2.6925 0.8325 ;
        RECT 2.5875 0.2175 2.6175 0.3825 ;
        RECT 2.5875 0.6675 2.6175 0.8325 ;
        END
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1125 0.2025 0.1425 0.3225 ;
        RECT 0.1125 0.6675 0.1425 0.8325 ;
        RECT 0.0375 0.2025 0.1125 0.8325 ;
        END
    END CO
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 2.2575 0.4050 2.3625 0.5550 ;
        RECT 1.6200 0.4800 2.2575 0.5550 ;
        RECT 1.5450 0.4800 1.6200 0.6375 ;
        RECT 0.8625 0.5625 1.5450 0.6375 ;
        VIA 2.3100 0.4800 VIA12_square ;
        VIA 1.6425 0.5175 VIA12_square ;
        VIA 0.9450 0.6000 VIA12_square ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.8550 0.4125 1.3200 0.4875 ;
        VIA 1.0950 0.4500 VIA12_square ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 2.4750 -0.0750 2.7300 0.0750 ;
        RECT 2.3700 -0.0750 2.4750 0.2250 ;
        RECT 1.4250 -0.0750 2.3700 0.0750 ;
        RECT 1.3050 -0.0750 1.4250 0.1800 ;
        RECT 0.9900 -0.0750 1.3050 0.0750 ;
        RECT 0.9000 -0.0750 0.9900 0.3000 ;
        RECT 0.3750 -0.0750 0.9000 0.0750 ;
        RECT 0.2550 -0.0750 0.3750 0.1875 ;
        RECT 0.0000 -0.0750 0.2550 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 2.4750 0.9750 2.7300 1.1250 ;
        RECT 2.3550 0.8700 2.4750 1.1250 ;
        RECT 1.2150 0.9750 2.3550 1.1250 ;
        RECT 1.0950 0.8700 1.2150 1.1250 ;
        RECT 0.7725 0.9750 1.0950 1.1250 ;
        RECT 0.6975 0.7500 0.7725 1.1250 ;
        RECT 0.3750 0.9750 0.6975 1.1250 ;
        RECT 0.2550 0.8700 0.3750 1.1250 ;
        RECT 0.0000 0.9750 0.2550 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 2.5950 0.2550 2.6550 0.3150 ;
        RECT 2.5950 0.7275 2.6550 0.7875 ;
        RECT 2.4825 0.4875 2.5425 0.5475 ;
        RECT 2.3850 0.1350 2.4450 0.1950 ;
        RECT 2.3850 0.8700 2.4450 0.9300 ;
        RECT 2.2725 0.4650 2.3325 0.5250 ;
        RECT 2.1750 0.1575 2.2350 0.2175 ;
        RECT 2.1750 0.7275 2.2350 0.7875 ;
        RECT 1.9650 0.2250 2.0250 0.2850 ;
        RECT 1.9650 0.8325 2.0250 0.8925 ;
        RECT 1.8600 0.4950 1.9200 0.5550 ;
        RECT 1.7550 0.1725 1.8150 0.2325 ;
        RECT 1.7550 0.6675 1.8150 0.7275 ;
        RECT 1.6500 0.4425 1.7100 0.5025 ;
        RECT 1.5450 0.6675 1.6050 0.7275 ;
        RECT 1.4325 0.4125 1.4925 0.4725 ;
        RECT 1.3350 0.1200 1.3950 0.1800 ;
        RECT 1.3350 0.8250 1.3950 0.8850 ;
        RECT 1.2300 0.4125 1.2900 0.4725 ;
        RECT 1.2300 0.6525 1.2900 0.7125 ;
        RECT 1.1250 0.2400 1.1850 0.3000 ;
        RECT 1.1250 0.8700 1.1850 0.9300 ;
        RECT 1.0200 0.4275 1.0800 0.4875 ;
        RECT 0.9150 0.1950 0.9750 0.2550 ;
        RECT 0.9150 0.7875 0.9750 0.8475 ;
        RECT 0.8100 0.4275 0.8700 0.4875 ;
        RECT 0.7050 0.2100 0.7650 0.2700 ;
        RECT 0.7050 0.7875 0.7650 0.8475 ;
        RECT 0.6075 0.4275 0.6675 0.4875 ;
        RECT 0.4950 0.7275 0.5550 0.7875 ;
        RECT 0.3900 0.4950 0.4500 0.5550 ;
        RECT 0.2850 0.1200 0.3450 0.1800 ;
        RECT 0.2850 0.8700 0.3450 0.9300 ;
        RECT 0.1875 0.4800 0.2475 0.5400 ;
        RECT 0.0750 0.2325 0.1350 0.2925 ;
        RECT 0.0750 0.7200 0.1350 0.7800 ;
        LAYER M1 ;
        RECT 2.5125 0.4575 2.5425 0.5775 ;
        RECT 2.4375 0.4575 2.5125 0.7950 ;
        RECT 2.3625 0.3000 2.4675 0.3825 ;
        RECT 2.3100 0.6900 2.4375 0.7950 ;
        RECT 2.2725 0.3000 2.3625 0.5850 ;
        RECT 2.1975 0.1500 2.2650 0.2250 ;
        RECT 2.1975 0.6675 2.2350 0.8175 ;
        RECT 2.1600 0.1500 2.1975 0.8175 ;
        RECT 2.1225 0.1500 2.1600 0.7425 ;
        RECT 1.8300 0.4950 2.1225 0.5700 ;
        RECT 1.4100 0.8250 2.0550 0.9000 ;
        RECT 1.9500 0.1800 2.0475 0.4200 ;
        RECT 1.7025 0.6450 2.0100 0.7500 ;
        RECT 1.8150 0.3300 1.9500 0.4200 ;
        RECT 1.5750 0.1500 1.8750 0.2550 ;
        RECT 1.7100 0.4650 1.7175 0.5700 ;
        RECT 1.5675 0.3300 1.7100 0.5700 ;
        RECT 1.5000 0.6450 1.6275 0.7500 ;
        RECT 1.4925 0.6450 1.5000 0.7200 ;
        RECT 1.4175 0.2550 1.4925 0.7200 ;
        RECT 1.2075 0.2550 1.4175 0.3375 ;
        RECT 1.2075 0.6450 1.4175 0.7200 ;
        RECT 1.3050 0.7950 1.4100 0.9000 ;
        RECT 1.2075 0.4125 1.3200 0.5175 ;
        RECT 1.1025 0.2100 1.2075 0.3375 ;
        RECT 0.5700 0.4125 1.2075 0.4875 ;
        RECT 1.1325 0.6450 1.2075 0.7950 ;
        RECT 0.9900 0.7200 1.1325 0.7950 ;
        RECT 0.4650 0.5625 1.0275 0.6375 ;
        RECT 0.9075 0.7200 0.9900 0.8775 ;
        RECT 0.6750 0.2025 0.7950 0.3375 ;
        RECT 0.3150 0.2625 0.6750 0.3375 ;
        RECT 0.3150 0.7200 0.5925 0.7950 ;
        RECT 0.3900 0.4650 0.4650 0.6375 ;
        RECT 0.2400 0.2625 0.3150 0.7950 ;
        RECT 0.1875 0.4500 0.2400 0.5700 ;
        LAYER VIA1 ;
        RECT 2.3550 0.7125 2.4300 0.7875 ;
        RECT 1.8975 0.3300 1.9725 0.4050 ;
        RECT 1.8825 0.6675 1.9575 0.7425 ;
        RECT 1.6800 0.1575 1.7550 0.2325 ;
        RECT 1.3725 0.2625 1.4475 0.3375 ;
        LAYER M2 ;
        RECT 1.9950 0.7125 2.5050 0.7875 ;
        RECT 1.5600 0.3300 2.0175 0.4050 ;
        RECT 1.8450 0.6525 1.9950 0.7875 ;
        RECT 0.7050 0.7125 1.8450 0.7875 ;
        RECT 1.6350 0.1125 1.8000 0.2475 ;
        RECT 0.7050 0.1125 1.6350 0.1875 ;
        RECT 1.4775 0.2625 1.5600 0.4050 ;
        RECT 1.3275 0.2625 1.4775 0.3375 ;
        RECT 0.6300 0.1125 0.7050 0.7875 ;
    END
END HA1_1010


MACRO IND2_0010
    CLASS CORE ;
    FOREIGN IND2_0010 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.2500 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 2.3625 0.2925 2.5200 0.4125 ;
        RECT 2.3625 0.6450 2.5200 0.7650 ;
        RECT 2.0475 0.2925 2.3625 0.7650 ;
        RECT 1.8900 0.2925 2.0475 0.4125 ;
        RECT 1.8900 0.6450 2.0475 0.7650 ;
        VIA 2.3625 0.3525 VIA12_slot ;
        VIA 2.3625 0.7050 VIA12_slot ;
        VIA 2.0475 0.3525 VIA12_slot ;
        VIA 2.0475 0.7050 VIA12_slot ;
        END
    END ZN
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 4.9125 0.4125 5.0775 0.6375 ;
        RECT 2.6700 0.4125 4.9125 0.5250 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1425 0.4500 0.6600 0.5700 ;
        RECT 0.0675 0.3675 0.1425 0.6825 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 4.9950 -0.0750 5.2500 0.0750 ;
        RECT 4.8750 -0.0750 4.9950 0.1875 ;
        RECT 4.5750 -0.0750 4.8750 0.0750 ;
        RECT 4.4550 -0.0750 4.5750 0.1875 ;
        RECT 4.1550 -0.0750 4.4550 0.0750 ;
        RECT 4.0350 -0.0750 4.1550 0.1875 ;
        RECT 3.7350 -0.0750 4.0350 0.0750 ;
        RECT 3.6150 -0.0750 3.7350 0.1875 ;
        RECT 3.3150 -0.0750 3.6150 0.0750 ;
        RECT 3.1950 -0.0750 3.3150 0.1875 ;
        RECT 2.8950 -0.0750 3.1950 0.0750 ;
        RECT 2.7750 -0.0750 2.8950 0.1875 ;
        RECT 0.5850 -0.0750 2.7750 0.0750 ;
        RECT 0.4650 -0.0750 0.5850 0.2250 ;
        RECT 0.1575 -0.0750 0.4650 0.0750 ;
        RECT 0.0525 -0.0750 0.1575 0.2625 ;
        RECT 0.0000 -0.0750 0.0525 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 5.1825 0.9750 5.2500 1.1250 ;
        RECT 5.1075 0.7800 5.1825 1.1250 ;
        RECT 4.7850 0.9750 5.1075 1.1250 ;
        RECT 4.6650 0.8625 4.7850 1.1250 ;
        RECT 4.3650 0.9750 4.6650 1.1250 ;
        RECT 4.2450 0.8625 4.3650 1.1250 ;
        RECT 3.9450 0.9750 4.2450 1.1250 ;
        RECT 3.8250 0.8625 3.9450 1.1250 ;
        RECT 3.5250 0.9750 3.8250 1.1250 ;
        RECT 3.4050 0.8625 3.5250 1.1250 ;
        RECT 3.1050 0.9750 3.4050 1.1250 ;
        RECT 2.9850 0.8625 3.1050 1.1250 ;
        RECT 2.6850 0.9750 2.9850 1.1250 ;
        RECT 2.5650 0.8625 2.6850 1.1250 ;
        RECT 2.2650 0.9750 2.5650 1.1250 ;
        RECT 2.1450 0.8625 2.2650 1.1250 ;
        RECT 1.8450 0.9750 2.1450 1.1250 ;
        RECT 1.7250 0.8625 1.8450 1.1250 ;
        RECT 1.4250 0.9750 1.7250 1.1250 ;
        RECT 1.3050 0.8625 1.4250 1.1250 ;
        RECT 0.9975 0.9750 1.3050 1.1250 ;
        RECT 0.8925 0.7875 0.9975 1.1250 ;
        RECT 0.5850 0.9750 0.8925 1.1250 ;
        RECT 0.4650 0.8250 0.5850 1.1250 ;
        RECT 0.1575 0.9750 0.4650 1.1250 ;
        RECT 0.0525 0.7875 0.1575 1.1250 ;
        RECT 0.0000 0.9750 0.0525 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 5.1150 0.2100 5.1750 0.2700 ;
        RECT 5.1150 0.8325 5.1750 0.8925 ;
        RECT 5.0100 0.4650 5.0700 0.5250 ;
        RECT 4.9050 0.1275 4.9650 0.1875 ;
        RECT 4.9050 0.8175 4.9650 0.8775 ;
        RECT 4.8000 0.4650 4.8600 0.5250 ;
        RECT 4.6950 0.2700 4.7550 0.3300 ;
        RECT 4.6950 0.8625 4.7550 0.9225 ;
        RECT 4.5900 0.4650 4.6500 0.5250 ;
        RECT 4.4850 0.1275 4.5450 0.1875 ;
        RECT 4.4850 0.8175 4.5450 0.8775 ;
        RECT 4.3800 0.4650 4.4400 0.5250 ;
        RECT 4.2750 0.2700 4.3350 0.3300 ;
        RECT 4.2750 0.8625 4.3350 0.9225 ;
        RECT 4.1700 0.4650 4.2300 0.5250 ;
        RECT 4.0650 0.1275 4.1250 0.1875 ;
        RECT 4.0650 0.8175 4.1250 0.8775 ;
        RECT 3.9600 0.4650 4.0200 0.5250 ;
        RECT 3.8550 0.2700 3.9150 0.3300 ;
        RECT 3.8550 0.8625 3.9150 0.9225 ;
        RECT 3.7500 0.4650 3.8100 0.5250 ;
        RECT 3.6450 0.1275 3.7050 0.1875 ;
        RECT 3.6450 0.8175 3.7050 0.8775 ;
        RECT 3.5400 0.4650 3.6000 0.5250 ;
        RECT 3.4350 0.2700 3.4950 0.3300 ;
        RECT 3.4350 0.8625 3.4950 0.9225 ;
        RECT 3.3300 0.4650 3.3900 0.5250 ;
        RECT 3.2250 0.1275 3.2850 0.1875 ;
        RECT 3.2250 0.6975 3.2850 0.7575 ;
        RECT 3.1200 0.4650 3.1800 0.5250 ;
        RECT 3.0150 0.2700 3.0750 0.3300 ;
        RECT 3.0150 0.8625 3.0750 0.9225 ;
        RECT 2.9100 0.4650 2.9700 0.5250 ;
        RECT 2.8050 0.1275 2.8650 0.1875 ;
        RECT 2.8050 0.6975 2.8650 0.7575 ;
        RECT 2.7000 0.4650 2.7600 0.5250 ;
        RECT 2.5950 0.1575 2.6550 0.2175 ;
        RECT 2.5950 0.8625 2.6550 0.9225 ;
        RECT 2.4900 0.4800 2.5500 0.5400 ;
        RECT 2.3850 0.3000 2.4450 0.3600 ;
        RECT 2.3850 0.6975 2.4450 0.7575 ;
        RECT 2.2800 0.4800 2.3400 0.5400 ;
        RECT 2.1750 0.1575 2.2350 0.2175 ;
        RECT 2.1750 0.8625 2.2350 0.9225 ;
        RECT 2.0700 0.4800 2.1300 0.5400 ;
        RECT 1.9650 0.3000 2.0250 0.3600 ;
        RECT 1.9650 0.6975 2.0250 0.7575 ;
        RECT 1.8600 0.4800 1.9200 0.5400 ;
        RECT 1.7550 0.1575 1.8150 0.2175 ;
        RECT 1.7550 0.8625 1.8150 0.9225 ;
        RECT 1.6500 0.4800 1.7100 0.5400 ;
        RECT 1.5450 0.3000 1.6050 0.3600 ;
        RECT 1.5450 0.6975 1.6050 0.7575 ;
        RECT 1.4400 0.4800 1.5000 0.5400 ;
        RECT 1.3350 0.1575 1.3950 0.2175 ;
        RECT 1.3350 0.8625 1.3950 0.9225 ;
        RECT 1.2300 0.4800 1.2900 0.5400 ;
        RECT 1.1250 0.3000 1.1850 0.3600 ;
        RECT 1.1250 0.6975 1.1850 0.7575 ;
        RECT 1.0200 0.4800 1.0800 0.5400 ;
        RECT 0.9150 0.1800 0.9750 0.2400 ;
        RECT 0.9150 0.8175 0.9750 0.8775 ;
        RECT 0.7050 0.3000 0.7650 0.3600 ;
        RECT 0.7050 0.6675 0.7650 0.7275 ;
        RECT 0.6000 0.4800 0.6600 0.5400 ;
        RECT 0.4950 0.1650 0.5550 0.2250 ;
        RECT 0.4950 0.8325 0.5550 0.8925 ;
        RECT 0.3900 0.4800 0.4500 0.5400 ;
        RECT 0.2850 0.2925 0.3450 0.3525 ;
        RECT 0.2850 0.6675 0.3450 0.7275 ;
        RECT 0.1800 0.4800 0.2400 0.5400 ;
        RECT 0.0750 0.1725 0.1350 0.2325 ;
        RECT 0.0750 0.8175 0.1350 0.8775 ;
        LAYER M1 ;
        RECT 5.1075 0.1800 5.1825 0.3375 ;
        RECT 2.6925 0.2625 5.1075 0.3375 ;
        RECT 4.8825 0.7125 4.9875 0.9000 ;
        RECT 4.8375 0.7125 4.8825 0.7875 ;
        RECT 4.5675 0.6675 4.8375 0.7875 ;
        RECT 4.4625 0.6675 4.5675 0.9000 ;
        RECT 4.1475 0.6675 4.4625 0.7875 ;
        RECT 4.0425 0.6675 4.1475 0.9000 ;
        RECT 3.7275 0.6675 4.0425 0.7875 ;
        RECT 3.6225 0.6675 3.7275 0.9000 ;
        RECT 1.1175 0.6675 3.6225 0.7875 ;
        RECT 2.6175 0.1500 2.6925 0.3375 ;
        RECT 0.9975 0.1500 2.6175 0.2250 ;
        RECT 0.8100 0.4800 2.5800 0.5850 ;
        RECT 1.0950 0.3000 2.5425 0.4050 ;
        RECT 0.8925 0.1500 0.9975 0.2700 ;
        RECT 0.7350 0.3000 0.8100 0.7500 ;
        RECT 0.3750 0.3000 0.7350 0.3750 ;
        RECT 0.2550 0.6450 0.7350 0.7500 ;
        RECT 0.2625 0.2700 0.3750 0.3750 ;
        LAYER M2 ;
        RECT 2.3925 0.2925 2.5200 0.4125 ;
        RECT 2.3925 0.6450 2.5200 0.7650 ;
        RECT 1.8900 0.2925 2.0175 0.4125 ;
        RECT 1.8900 0.6450 2.0175 0.7650 ;
    END
END IND2_0010


MACRO IND2_0011
    CLASS CORE ;
    FOREIGN IND2_0011 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.2600 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 0.9075 0.1125 0.9975 0.1875 ;
        RECT 0.8325 0.1125 0.9075 0.9375 ;
        RECT 0.3675 0.8625 0.8325 0.9375 ;
        VIA 0.8700 0.2025 VIA12_square ;
        VIA 0.8700 0.6900 VIA12_square ;
        END
    END ZN
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.6825 0.1125 0.7575 0.6900 ;
        RECT 0.2175 0.1125 0.6825 0.1875 ;
        VIA 0.7200 0.5100 VIA12_square ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.0975 0.5625 0.5625 0.6375 ;
        VIA 0.1800 0.6000 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.2000 -0.0750 1.2600 0.0750 ;
        RECT 1.1250 -0.0750 1.2000 0.2475 ;
        RECT 0.3750 -0.0750 1.1250 0.0750 ;
        RECT 0.2550 -0.0750 0.3750 0.1875 ;
        RECT 0.0000 -0.0750 0.2550 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.2075 0.9750 1.2600 1.1250 ;
        RECT 1.1025 0.8100 1.2075 1.1250 ;
        RECT 0.7950 0.9750 1.1025 1.1250 ;
        RECT 0.6750 0.8325 0.7950 1.1250 ;
        RECT 0.3750 0.9750 0.6750 1.1250 ;
        RECT 0.2550 0.8625 0.3750 1.1250 ;
        RECT 0.0000 0.9750 0.2550 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.1250 0.1575 1.1850 0.2175 ;
        RECT 1.1250 0.8325 1.1850 0.8925 ;
        RECT 1.0200 0.4800 1.0800 0.5400 ;
        RECT 0.9150 0.7425 0.9750 0.8025 ;
        RECT 0.8100 0.4950 0.8700 0.5550 ;
        RECT 0.7050 0.1725 0.7650 0.2325 ;
        RECT 0.7050 0.8400 0.7650 0.9000 ;
        RECT 0.6000 0.4950 0.6600 0.5550 ;
        RECT 0.4950 0.7425 0.5550 0.8025 ;
        RECT 0.3900 0.4800 0.4500 0.5400 ;
        RECT 0.2850 0.1275 0.3450 0.1875 ;
        RECT 0.2850 0.8625 0.3450 0.9225 ;
        RECT 0.1800 0.4800 0.2400 0.5400 ;
        RECT 0.0750 0.2475 0.1350 0.3075 ;
        RECT 0.0750 0.7425 0.1350 0.8025 ;
        LAYER M1 ;
        RECT 1.0425 0.4575 1.1025 0.5625 ;
        RECT 0.9675 0.3225 1.0425 0.5625 ;
        RECT 0.6750 0.1500 1.0200 0.2475 ;
        RECT 0.9075 0.6525 0.9825 0.8325 ;
        RECT 0.4500 0.3225 0.9675 0.3975 ;
        RECT 0.5625 0.6525 0.9075 0.7275 ;
        RECT 0.5775 0.4725 0.8925 0.5775 ;
        RECT 0.4875 0.6525 0.5625 0.8325 ;
        RECT 0.4125 0.3225 0.4500 0.5700 ;
        RECT 0.3375 0.2625 0.4125 0.7875 ;
        RECT 0.1425 0.2625 0.3375 0.3375 ;
        RECT 0.1425 0.7125 0.3375 0.7875 ;
        RECT 0.0975 0.4125 0.2625 0.6375 ;
        RECT 0.0675 0.2175 0.1425 0.3375 ;
        RECT 0.0675 0.7125 0.1425 0.8325 ;
    END
END IND2_0011


MACRO IND2_0111
    CLASS CORE ;
    FOREIGN IND2_0111 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.1000 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 1.2075 0.2625 1.5225 0.7350 ;
        VIA 1.3650 0.3450 VIA12_slot ;
        VIA 1.3650 0.6525 VIA12_slot ;
        END
    END ZN
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.9825 0.2625 1.0575 0.6075 ;
        RECT 0.5625 0.2625 0.9825 0.3375 ;
        VIA 1.0200 0.5025 VIA12_square ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.0975 0.5625 0.5625 0.6375 ;
        VIA 0.1800 0.6000 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 2.0325 -0.0750 2.1000 0.0750 ;
        RECT 1.9575 -0.0750 2.0325 0.2625 ;
        RECT 0.7950 -0.0750 1.9575 0.0750 ;
        RECT 0.6750 -0.0750 0.7950 0.1800 ;
        RECT 0.3750 -0.0750 0.6750 0.0750 ;
        RECT 0.2550 -0.0750 0.3750 0.1950 ;
        RECT 0.0000 -0.0750 0.2550 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 2.0475 0.9750 2.1000 1.1250 ;
        RECT 1.9425 0.6450 2.0475 1.1250 ;
        RECT 1.6275 0.9750 1.9425 1.1250 ;
        RECT 1.5225 0.8100 1.6275 1.1250 ;
        RECT 1.2075 0.9750 1.5225 1.1250 ;
        RECT 1.1025 0.8100 1.2075 1.1250 ;
        RECT 0.7875 0.9750 1.1025 1.1250 ;
        RECT 0.6825 0.8100 0.7875 1.1250 ;
        RECT 0.3750 0.9750 0.6825 1.1250 ;
        RECT 0.2550 0.8700 0.3750 1.1250 ;
        RECT 0.0000 0.9750 0.2550 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.9650 0.1725 2.0250 0.2325 ;
        RECT 1.9650 0.6675 2.0250 0.7275 ;
        RECT 1.9650 0.8325 2.0250 0.8925 ;
        RECT 1.8600 0.4650 1.9200 0.5250 ;
        RECT 1.7550 0.1575 1.8150 0.2175 ;
        RECT 1.7550 0.6525 1.8150 0.7125 ;
        RECT 1.6500 0.4725 1.7100 0.5325 ;
        RECT 1.5450 0.3000 1.6050 0.3600 ;
        RECT 1.5450 0.8325 1.6050 0.8925 ;
        RECT 1.4400 0.4725 1.5000 0.5325 ;
        RECT 1.3350 0.1575 1.3950 0.2175 ;
        RECT 1.3350 0.6450 1.3950 0.7050 ;
        RECT 1.2300 0.4725 1.2900 0.5325 ;
        RECT 1.1250 0.3000 1.1850 0.3600 ;
        RECT 1.1250 0.8325 1.1850 0.8925 ;
        RECT 1.0200 0.4725 1.0800 0.5325 ;
        RECT 0.9150 0.2250 0.9750 0.2850 ;
        RECT 0.9150 0.6450 0.9750 0.7050 ;
        RECT 0.8025 0.4650 0.8625 0.5250 ;
        RECT 0.7050 0.1200 0.7650 0.1800 ;
        RECT 0.7050 0.8325 0.7650 0.8925 ;
        RECT 0.6000 0.4650 0.6600 0.5250 ;
        RECT 0.4950 0.2400 0.5550 0.3000 ;
        RECT 0.4950 0.7275 0.5550 0.7875 ;
        RECT 0.3900 0.4650 0.4500 0.5250 ;
        RECT 0.2850 0.1350 0.3450 0.1950 ;
        RECT 0.2850 0.8700 0.3450 0.9300 ;
        RECT 0.1800 0.4800 0.2400 0.5400 ;
        RECT 0.0750 0.2550 0.1350 0.3150 ;
        RECT 0.0750 0.7500 0.1350 0.8100 ;
        LAYER M1 ;
        RECT 1.8450 0.3900 2.0400 0.5550 ;
        RECT 0.9825 0.1500 1.8450 0.2250 ;
        RECT 1.7325 0.6300 1.8375 0.7350 ;
        RECT 1.0275 0.4650 1.7400 0.5400 ;
        RECT 1.0950 0.3000 1.7325 0.3900 ;
        RECT 0.9150 0.6150 1.7325 0.7350 ;
        RECT 0.9375 0.4350 1.0275 0.5400 ;
        RECT 0.9075 0.1500 0.9825 0.3300 ;
        RECT 0.5625 0.6300 0.9150 0.7350 ;
        RECT 0.5625 0.2550 0.9075 0.3300 ;
        RECT 0.4125 0.4350 0.8625 0.5550 ;
        RECT 0.4875 0.2100 0.5625 0.3300 ;
        RECT 0.4875 0.6300 0.5625 0.8250 ;
        RECT 0.3375 0.2700 0.4125 0.7950 ;
        RECT 0.1425 0.2700 0.3375 0.3450 ;
        RECT 0.1425 0.7200 0.3375 0.7950 ;
        RECT 0.0975 0.4200 0.2625 0.6450 ;
        RECT 0.0675 0.2250 0.1425 0.3450 ;
        RECT 0.0675 0.7200 0.1425 0.8400 ;
        LAYER VIA1 ;
        RECT 1.8900 0.4125 1.9650 0.4875 ;
        RECT 0.7125 0.4575 0.7875 0.5325 ;
        LAYER M2 ;
        RECT 1.7475 0.4125 2.0100 0.4875 ;
        RECT 1.6725 0.4125 1.7475 0.9375 ;
        RECT 0.7725 0.8625 1.6725 0.9375 ;
        RECT 0.7725 0.4125 0.8025 0.5775 ;
        RECT 0.6975 0.4125 0.7725 0.9375 ;
    END
END IND2_0111


MACRO IND2_1000
    CLASS CORE ;
    FOREIGN IND2_1000 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.8400 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.7275 0.1500 0.8025 0.7425 ;
        RECT 0.6750 0.1500 0.7275 0.2625 ;
        RECT 0.5625 0.6675 0.7275 0.7425 ;
        RECT 0.4875 0.6675 0.5625 0.8700 ;
        END
    END ZN
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.5625 0.3375 0.6525 0.5925 ;
        RECT 0.5475 0.2175 0.5625 0.5925 ;
        RECT 0.4875 0.2175 0.5475 0.4125 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.0975 0.5625 0.5625 0.6375 ;
        VIA 0.1800 0.6000 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.3750 -0.0750 0.8400 0.0750 ;
        RECT 0.2550 -0.0750 0.3750 0.2175 ;
        RECT 0.0000 -0.0750 0.2550 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.7950 0.9750 0.8400 1.1250 ;
        RECT 0.6750 0.8175 0.7950 1.1250 ;
        RECT 0.3750 0.9750 0.6750 1.1250 ;
        RECT 0.2550 0.8625 0.3750 1.1250 ;
        RECT 0.0000 0.9750 0.2550 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 0.7050 0.1575 0.7650 0.2175 ;
        RECT 0.7050 0.8325 0.7650 0.8925 ;
        RECT 0.5925 0.4950 0.6525 0.5550 ;
        RECT 0.4950 0.7800 0.5550 0.8400 ;
        RECT 0.3825 0.5025 0.4425 0.5625 ;
        RECT 0.2850 0.1500 0.3450 0.2100 ;
        RECT 0.2850 0.8700 0.3450 0.9300 ;
        RECT 0.1800 0.4800 0.2400 0.5400 ;
        RECT 0.0750 0.1575 0.1350 0.2175 ;
        RECT 0.0750 0.8175 0.1350 0.8775 ;
        LAYER M1 ;
        RECT 0.4125 0.4725 0.4425 0.5925 ;
        RECT 0.3375 0.2925 0.4125 0.7875 ;
        RECT 0.1650 0.2925 0.3375 0.3675 ;
        RECT 0.1575 0.7125 0.3375 0.7875 ;
        RECT 0.0975 0.4425 0.2625 0.6375 ;
        RECT 0.0450 0.1500 0.1650 0.3675 ;
        RECT 0.0525 0.7125 0.1575 0.9000 ;
    END
END IND2_1000


MACRO IND2_1010
    CLASS CORE ;
    FOREIGN IND2_1010 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.8400 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.7275 0.1650 0.8025 0.7425 ;
        RECT 0.6975 0.1650 0.7275 0.2850 ;
        RECT 0.5625 0.6675 0.7275 0.7425 ;
        RECT 0.4875 0.6675 0.5625 0.8325 ;
        END
    END ZN
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.6225 0.4575 0.6525 0.5925 ;
        RECT 0.5475 0.2175 0.6225 0.5925 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.2625 0.2625 0.3825 0.3975 ;
        RECT 0.2175 0.2625 0.2625 0.5775 ;
        RECT 0.1875 0.3375 0.2175 0.5775 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.3750 -0.0750 0.8400 0.0750 ;
        RECT 0.2550 -0.0750 0.3750 0.1875 ;
        RECT 0.0000 -0.0750 0.2550 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.7950 0.9750 0.8400 1.1250 ;
        RECT 0.6750 0.8175 0.7950 1.1250 ;
        RECT 0.3750 0.9750 0.6750 1.1250 ;
        RECT 0.2550 0.8625 0.3750 1.1250 ;
        RECT 0.0000 0.9750 0.2550 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 0.7050 0.1950 0.7650 0.2550 ;
        RECT 0.7050 0.8325 0.7650 0.8925 ;
        RECT 0.5925 0.4950 0.6525 0.5550 ;
        RECT 0.4950 0.7425 0.5550 0.8025 ;
        RECT 0.3825 0.5025 0.4425 0.5625 ;
        RECT 0.2850 0.1200 0.3450 0.1800 ;
        RECT 0.2850 0.8700 0.3450 0.9300 ;
        RECT 0.1875 0.4800 0.2475 0.5400 ;
        RECT 0.0750 0.1800 0.1350 0.2400 ;
        RECT 0.0750 0.7200 0.1350 0.7800 ;
        LAYER M1 ;
        RECT 0.4125 0.4725 0.4425 0.5925 ;
        RECT 0.3375 0.4725 0.4125 0.7875 ;
        RECT 0.1125 0.7125 0.3375 0.7875 ;
        RECT 0.1125 0.1500 0.1425 0.2700 ;
        RECT 0.0375 0.1500 0.1125 0.7875 ;
    END
END IND2_1010


MACRO IND3_0011
    CLASS CORE ;
    FOREIGN IND3_0011 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.8900 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 0.2175 0.7125 0.7725 0.7875 ;
        VIA 0.5250 0.7500 VIA12_square ;
        END
    END ZN
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.1025 0.4425 1.2075 0.6375 ;
        RECT 0.6525 0.5625 1.1025 0.6375 ;
        VIA 1.1550 0.5250 VIA12_square ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.4325 0.4650 1.5375 0.7875 ;
        RECT 0.9975 0.7125 1.4325 0.7875 ;
        VIA 1.4850 0.5475 VIA12_square ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.0900 0.4125 0.5550 0.4875 ;
        VIA 0.1725 0.4500 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.7800 -0.0750 1.8900 0.0750 ;
        RECT 0.6750 -0.0750 0.7800 0.2475 ;
        RECT 0.3750 -0.0750 0.6750 0.0750 ;
        RECT 0.2550 -0.0750 0.3750 0.1875 ;
        RECT 0.0000 -0.0750 0.2550 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.8375 0.9750 1.8900 1.1250 ;
        RECT 1.7325 0.8100 1.8375 1.1250 ;
        RECT 1.4250 0.9750 1.7325 1.1250 ;
        RECT 1.3050 0.8250 1.4250 1.1250 ;
        RECT 1.0050 0.9750 1.3050 1.1250 ;
        RECT 0.8850 0.8250 1.0050 1.1250 ;
        RECT 0.7950 0.9750 0.8850 1.1250 ;
        RECT 0.6750 0.8250 0.7950 1.1250 ;
        RECT 0.3750 0.9750 0.6750 1.1250 ;
        RECT 0.2550 0.8550 0.3750 1.1250 ;
        RECT 0.0000 0.9750 0.2550 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.7550 0.1725 1.8150 0.2325 ;
        RECT 1.7550 0.8325 1.8150 0.8925 ;
        RECT 1.6500 0.4950 1.7100 0.5550 ;
        RECT 1.5450 0.3150 1.6050 0.3750 ;
        RECT 1.5450 0.7125 1.6050 0.7725 ;
        RECT 1.4400 0.4950 1.5000 0.5550 ;
        RECT 1.3350 0.1575 1.3950 0.2175 ;
        RECT 1.3350 0.8325 1.3950 0.8925 ;
        RECT 1.2300 0.4950 1.2900 0.5550 ;
        RECT 1.1250 0.3075 1.1850 0.3675 ;
        RECT 1.1250 0.7125 1.1850 0.7725 ;
        RECT 1.0200 0.4950 1.0800 0.5550 ;
        RECT 0.9150 0.1575 0.9750 0.2175 ;
        RECT 0.9150 0.8325 0.9750 0.8925 ;
        RECT 0.7050 0.1575 0.7650 0.2175 ;
        RECT 0.7050 0.8325 0.7650 0.8925 ;
        RECT 0.6000 0.4950 0.6600 0.5550 ;
        RECT 0.4950 0.2925 0.5550 0.3525 ;
        RECT 0.4950 0.7125 0.5550 0.7725 ;
        RECT 0.3900 0.4950 0.4500 0.5550 ;
        RECT 0.2850 0.1275 0.3450 0.1875 ;
        RECT 0.2850 0.8550 0.3450 0.9150 ;
        RECT 0.1800 0.4800 0.2400 0.5400 ;
        RECT 0.0750 0.2475 0.1350 0.3075 ;
        RECT 0.0750 0.7350 0.1350 0.7950 ;
        LAYER M1 ;
        RECT 1.7325 0.1500 1.8375 0.2550 ;
        RECT 1.3875 0.4800 1.7475 0.5850 ;
        RECT 0.8850 0.1500 1.7325 0.2250 ;
        RECT 1.4250 0.3000 1.6725 0.4050 ;
        RECT 1.5375 0.6600 1.6125 0.8325 ;
        RECT 1.1925 0.6600 1.5375 0.7350 ;
        RECT 1.3200 0.3000 1.4250 0.3900 ;
        RECT 0.9975 0.4725 1.3125 0.5775 ;
        RECT 0.9225 0.3000 1.2150 0.3750 ;
        RECT 1.1175 0.6600 1.1925 0.8325 ;
        RECT 0.9225 0.6600 1.1175 0.7350 ;
        RECT 0.8400 0.3000 0.9225 0.7350 ;
        RECT 0.5625 0.6600 0.8400 0.7350 ;
        RECT 0.6000 0.3225 0.7350 0.3975 ;
        RECT 0.4050 0.4875 0.6900 0.5625 ;
        RECT 0.4875 0.1500 0.6000 0.3975 ;
        RECT 0.4875 0.6600 0.5625 0.8325 ;
        RECT 0.3300 0.2625 0.4050 0.7800 ;
        RECT 0.1425 0.2625 0.3300 0.3375 ;
        RECT 0.1425 0.7050 0.3300 0.7800 ;
        RECT 0.0900 0.4125 0.2550 0.6300 ;
        RECT 0.0675 0.2175 0.1425 0.3375 ;
        RECT 0.0675 0.7050 0.1425 0.8250 ;
        LAYER VIA1 ;
        RECT 1.3725 0.3000 1.4475 0.3750 ;
        RECT 0.5100 0.2625 0.5850 0.3375 ;
        LAYER M2 ;
        RECT 1.3800 0.3000 1.4925 0.3750 ;
        RECT 1.3050 0.2625 1.3800 0.3750 ;
        RECT 0.4425 0.2625 1.3050 0.3375 ;
    END
END IND3_0011


MACRO IND3_0111
    CLASS CORE ;
    FOREIGN IND3_0111 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.1500 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 2.4675 0.2625 2.7825 0.7800 ;
        VIA 2.6250 0.3450 VIA12_slot ;
        VIA 2.6250 0.6975 VIA12_slot ;
        END
    END ZN
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 3.0075 0.3675 3.0825 0.6825 ;
        RECT 2.2575 0.4650 3.0075 0.5700 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.7475 0.4125 1.8225 0.5850 ;
        RECT 1.2825 0.4125 1.7475 0.4875 ;
        VIA 1.7850 0.5025 VIA12_square ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.0900 0.4125 0.5550 0.4875 ;
        VIA 0.1725 0.4500 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.2000 -0.0750 3.1500 0.0750 ;
        RECT 1.0950 -0.0750 1.2000 0.2475 ;
        RECT 0.7875 -0.0750 1.0950 0.0750 ;
        RECT 0.6825 -0.0750 0.7875 0.2400 ;
        RECT 0.3750 -0.0750 0.6825 0.0750 ;
        RECT 0.2550 -0.0750 0.3750 0.1875 ;
        RECT 0.0000 -0.0750 0.2550 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 3.0825 0.9750 3.1500 1.1250 ;
        RECT 3.0075 0.7875 3.0825 1.1250 ;
        RECT 2.6850 0.9750 3.0075 1.1250 ;
        RECT 2.5650 0.8250 2.6850 1.1250 ;
        RECT 2.2650 0.9750 2.5650 1.1250 ;
        RECT 2.1450 0.8250 2.2650 1.1250 ;
        RECT 1.8450 0.9750 2.1450 1.1250 ;
        RECT 1.7250 0.8250 1.8450 1.1250 ;
        RECT 1.4250 0.9750 1.7250 1.1250 ;
        RECT 1.3050 0.8250 1.4250 1.1250 ;
        RECT 1.2150 0.9750 1.3050 1.1250 ;
        RECT 1.0950 0.8250 1.2150 1.1250 ;
        RECT 0.7950 0.9750 1.0950 1.1250 ;
        RECT 0.6750 0.8250 0.7950 1.1250 ;
        RECT 0.3750 0.9750 0.6750 1.1250 ;
        RECT 0.2550 0.8550 0.3750 1.1250 ;
        RECT 0.0000 0.9750 0.2550 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 3.0150 0.1725 3.0750 0.2325 ;
        RECT 3.0150 0.8175 3.0750 0.8775 ;
        RECT 2.9100 0.4875 2.9700 0.5475 ;
        RECT 2.8050 0.3150 2.8650 0.3750 ;
        RECT 2.8050 0.6675 2.8650 0.7275 ;
        RECT 2.7000 0.4875 2.7600 0.5475 ;
        RECT 2.5950 0.1575 2.6550 0.2175 ;
        RECT 2.5950 0.8325 2.6550 0.8925 ;
        RECT 2.4900 0.4875 2.5500 0.5475 ;
        RECT 2.3850 0.3150 2.4450 0.3750 ;
        RECT 2.3850 0.6675 2.4450 0.7275 ;
        RECT 2.2800 0.4875 2.3400 0.5475 ;
        RECT 2.1750 0.1575 2.2350 0.2175 ;
        RECT 2.1750 0.8325 2.2350 0.8925 ;
        RECT 2.0700 0.4875 2.1300 0.5475 ;
        RECT 1.9650 0.3075 2.0250 0.3675 ;
        RECT 1.9650 0.6675 2.0250 0.7275 ;
        RECT 1.8600 0.4875 1.9200 0.5475 ;
        RECT 1.7550 0.1575 1.8150 0.2175 ;
        RECT 1.7550 0.8325 1.8150 0.8925 ;
        RECT 1.6500 0.4875 1.7100 0.5475 ;
        RECT 1.5450 0.3075 1.6050 0.3675 ;
        RECT 1.5450 0.6675 1.6050 0.7275 ;
        RECT 1.4400 0.4875 1.5000 0.5475 ;
        RECT 1.3350 0.1575 1.3950 0.2175 ;
        RECT 1.3350 0.8325 1.3950 0.8925 ;
        RECT 1.1250 0.1575 1.1850 0.2175 ;
        RECT 1.1250 0.8325 1.1850 0.8925 ;
        RECT 1.0200 0.4950 1.0800 0.5550 ;
        RECT 0.9150 0.3225 0.9750 0.3825 ;
        RECT 0.9150 0.6675 0.9750 0.7275 ;
        RECT 0.8100 0.4950 0.8700 0.5550 ;
        RECT 0.7050 0.1575 0.7650 0.2175 ;
        RECT 0.7050 0.8325 0.7650 0.8925 ;
        RECT 0.6000 0.4950 0.6600 0.5550 ;
        RECT 0.4950 0.2925 0.5550 0.3525 ;
        RECT 0.4950 0.6900 0.5550 0.7500 ;
        RECT 0.3900 0.4950 0.4500 0.5550 ;
        RECT 0.2850 0.1275 0.3450 0.1875 ;
        RECT 0.2850 0.8550 0.3450 0.9150 ;
        RECT 0.1800 0.4800 0.2400 0.5400 ;
        RECT 0.0750 0.2475 0.1350 0.3075 ;
        RECT 0.0750 0.7350 0.1350 0.7950 ;
        LAYER M1 ;
        RECT 2.9925 0.1500 3.0975 0.2550 ;
        RECT 1.3050 0.1500 2.9925 0.2250 ;
        RECT 2.3550 0.3000 2.8950 0.3900 ;
        RECT 0.5625 0.6450 2.8875 0.7500 ;
        RECT 1.4175 0.4650 2.1525 0.5700 ;
        RECT 1.3425 0.3000 2.0550 0.3750 ;
        RECT 1.2600 0.3000 1.3425 0.3975 ;
        RECT 0.5625 0.3225 1.2600 0.3975 ;
        RECT 0.4050 0.4875 1.1100 0.5625 ;
        RECT 0.4875 0.2625 0.5625 0.3975 ;
        RECT 0.4875 0.6450 0.5625 0.7875 ;
        RECT 0.3300 0.2625 0.4050 0.7800 ;
        RECT 0.1425 0.2625 0.3300 0.3375 ;
        RECT 0.1425 0.7050 0.3300 0.7800 ;
        RECT 0.0900 0.4125 0.2550 0.6300 ;
        RECT 0.0675 0.2175 0.1425 0.3375 ;
        RECT 0.0675 0.7050 0.1425 0.8250 ;
    END
END IND3_0111


MACRO IND3_1000
    CLASS CORE ;
    FOREIGN IND3_1000 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.0500 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.9375 0.1500 1.0125 0.9000 ;
        RECT 0.9075 0.1500 0.9375 0.3825 ;
        RECT 0.9075 0.6675 0.9375 0.9000 ;
        RECT 0.5625 0.6675 0.9075 0.7425 ;
        RECT 0.4875 0.6675 0.5625 0.8700 ;
        END
    END ZN
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.4350 0.4125 0.9000 0.4875 ;
        VIA 0.7800 0.4500 VIA12_square ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.6225 0.1125 0.8400 0.1875 ;
        RECT 0.5175 0.1125 0.6225 0.2925 ;
        RECT 0.2700 0.1125 0.5175 0.1875 ;
        VIA 0.5700 0.2100 VIA12_square ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.0900 0.5625 0.5550 0.6375 ;
        VIA 0.1725 0.6000 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.3750 -0.0750 1.0500 0.0750 ;
        RECT 0.2550 -0.0750 0.3750 0.2025 ;
        RECT 0.0000 -0.0750 0.2550 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.7875 0.9750 1.0500 1.1250 ;
        RECT 0.6825 0.8175 0.7875 1.1250 ;
        RECT 0.3750 0.9750 0.6825 1.1250 ;
        RECT 0.2550 0.8625 0.3750 1.1250 ;
        RECT 0.0000 0.9750 0.2550 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 0.9150 0.1800 0.9750 0.2400 ;
        RECT 0.9150 0.8100 0.9750 0.8700 ;
        RECT 0.8025 0.4725 0.8625 0.5325 ;
        RECT 0.7050 0.8475 0.7650 0.9075 ;
        RECT 0.6000 0.4650 0.6600 0.5250 ;
        RECT 0.4950 0.7800 0.5550 0.8400 ;
        RECT 0.3900 0.4800 0.4500 0.5400 ;
        RECT 0.2850 0.1275 0.3450 0.1875 ;
        RECT 0.2850 0.8700 0.3450 0.9300 ;
        RECT 0.1800 0.4800 0.2400 0.5400 ;
        RECT 0.0750 0.1725 0.1350 0.2325 ;
        RECT 0.0750 0.8175 0.1350 0.8775 ;
        LAYER M1 ;
        RECT 0.8325 0.4425 0.8625 0.5925 ;
        RECT 0.7425 0.2775 0.8325 0.5925 ;
        RECT 0.5775 0.1725 0.6675 0.5625 ;
        RECT 0.4875 0.1725 0.5775 0.2775 ;
        RECT 0.4125 0.4575 0.4725 0.5625 ;
        RECT 0.3375 0.2775 0.4125 0.7875 ;
        RECT 0.1575 0.2775 0.3375 0.3525 ;
        RECT 0.1575 0.7125 0.3375 0.7875 ;
        RECT 0.0900 0.4275 0.2550 0.6375 ;
        RECT 0.0525 0.1500 0.1575 0.3525 ;
        RECT 0.0525 0.7125 0.1575 0.9000 ;
    END
END IND3_1000


MACRO IND3_1010
    CLASS CORE ;
    FOREIGN IND3_1010 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.0500 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.9375 0.2175 1.0125 0.8325 ;
        RECT 0.9075 0.2175 0.9375 0.3825 ;
        RECT 0.9075 0.6675 0.9375 0.8325 ;
        RECT 0.5625 0.6675 0.9075 0.7425 ;
        RECT 0.4875 0.6675 0.5625 0.8175 ;
        END
    END ZN
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.4350 0.4125 0.9000 0.4875 ;
        VIA 0.7800 0.4500 VIA12_square ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.6225 0.1125 0.8400 0.1875 ;
        RECT 0.5175 0.1125 0.6225 0.2925 ;
        RECT 0.2700 0.1125 0.5175 0.1875 ;
        VIA 0.5700 0.2100 VIA12_square ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.0900 0.5625 0.5550 0.6375 ;
        VIA 0.1725 0.6000 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.3750 -0.0750 1.0500 0.0750 ;
        RECT 0.2550 -0.0750 0.3750 0.2025 ;
        RECT 0.0000 -0.0750 0.2550 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.7875 0.9750 1.0500 1.1250 ;
        RECT 0.6825 0.8175 0.7875 1.1250 ;
        RECT 0.3750 0.9750 0.6825 1.1250 ;
        RECT 0.2550 0.8625 0.3750 1.1250 ;
        RECT 0.0000 0.9750 0.2550 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 0.9150 0.2700 0.9750 0.3300 ;
        RECT 0.9150 0.7200 0.9750 0.7800 ;
        RECT 0.8025 0.4725 0.8625 0.5325 ;
        RECT 0.7050 0.8475 0.7650 0.9075 ;
        RECT 0.6000 0.4650 0.6600 0.5250 ;
        RECT 0.4950 0.7125 0.5550 0.7725 ;
        RECT 0.3900 0.4800 0.4500 0.5400 ;
        RECT 0.2850 0.1275 0.3450 0.1875 ;
        RECT 0.2850 0.8700 0.3450 0.9300 ;
        RECT 0.1800 0.4800 0.2400 0.5400 ;
        RECT 0.0750 0.2625 0.1350 0.3225 ;
        RECT 0.0750 0.7500 0.1350 0.8100 ;
        LAYER M1 ;
        RECT 0.8325 0.4425 0.8625 0.5925 ;
        RECT 0.7425 0.2775 0.8325 0.5925 ;
        RECT 0.5775 0.1725 0.6675 0.5625 ;
        RECT 0.4875 0.1725 0.5775 0.2775 ;
        RECT 0.4125 0.4575 0.4725 0.5625 ;
        RECT 0.3375 0.2775 0.4125 0.7875 ;
        RECT 0.1425 0.2775 0.3375 0.3525 ;
        RECT 0.1425 0.7125 0.3375 0.7875 ;
        RECT 0.0900 0.4275 0.2550 0.6375 ;
        RECT 0.0675 0.2325 0.1425 0.3525 ;
        RECT 0.0675 0.7125 0.1425 0.8400 ;
    END
END IND3_1010


MACRO IND4_0011
    CLASS CORE ;
    FOREIGN IND4_0011 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.5200 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 2.3775 0.2100 2.4525 0.3750 ;
        RECT 1.9950 0.3000 2.3775 0.3750 ;
        RECT 2.1600 0.6450 2.2350 0.8325 ;
        RECT 1.9950 0.6450 2.1600 0.7200 ;
        RECT 1.9200 0.3000 1.9950 0.7200 ;
        RECT 1.6125 0.6450 1.9200 0.7200 ;
        RECT 1.5375 0.6450 1.6125 0.8325 ;
        RECT 1.1925 0.6450 1.5375 0.7200 ;
        RECT 1.1175 0.6450 1.1925 0.8325 ;
        RECT 0.5625 0.6450 1.1175 0.7200 ;
        RECT 0.4875 0.6450 0.5625 0.8325 ;
        END
    END ZN
    PIN B3
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.8600 0.5625 2.4300 0.6375 ;
        VIA 2.3475 0.6000 VIA12_square ;
        END
    END B3
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.5375 0.2625 1.6125 0.6075 ;
        RECT 1.0725 0.2625 1.5375 0.3375 ;
        VIA 1.5750 0.5250 VIA12_square ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.1175 0.4125 1.1925 0.6000 ;
        RECT 0.6525 0.4125 1.1175 0.4875 ;
        VIA 1.1550 0.5175 VIA12_square ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.0900 0.5625 0.5550 0.6375 ;
        VIA 0.1725 0.6000 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.7800 -0.0750 2.5200 0.0750 ;
        RECT 0.6750 -0.0750 0.7800 0.2475 ;
        RECT 0.3750 -0.0750 0.6750 0.0750 ;
        RECT 0.2550 -0.0750 0.3750 0.1950 ;
        RECT 0.0000 -0.0750 0.2550 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 2.4525 0.9750 2.5200 1.1250 ;
        RECT 2.3775 0.7875 2.4525 1.1250 ;
        RECT 2.0550 0.9750 2.3775 1.1250 ;
        RECT 1.9350 0.8250 2.0550 1.1250 ;
        RECT 1.8450 0.9750 1.9350 1.1250 ;
        RECT 1.7250 0.8250 1.8450 1.1250 ;
        RECT 1.4250 0.9750 1.7250 1.1250 ;
        RECT 1.3050 0.8250 1.4250 1.1250 ;
        RECT 1.0050 0.9750 1.3050 1.1250 ;
        RECT 0.8850 0.8250 1.0050 1.1250 ;
        RECT 0.7950 0.9750 0.8850 1.1250 ;
        RECT 0.6750 0.8250 0.7950 1.1250 ;
        RECT 0.3750 0.9750 0.6750 1.1250 ;
        RECT 0.2550 0.8625 0.3750 1.1250 ;
        RECT 0.0000 0.9750 0.2550 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 2.3850 0.2400 2.4450 0.3000 ;
        RECT 2.3850 0.8175 2.4450 0.8775 ;
        RECT 2.2800 0.4800 2.3400 0.5400 ;
        RECT 2.1750 0.1575 2.2350 0.2175 ;
        RECT 2.1750 0.7425 2.2350 0.8025 ;
        RECT 2.0700 0.4800 2.1300 0.5400 ;
        RECT 1.9650 0.3000 2.0250 0.3600 ;
        RECT 1.9650 0.8325 2.0250 0.8925 ;
        RECT 1.7550 0.3075 1.8150 0.3675 ;
        RECT 1.7550 0.8325 1.8150 0.8925 ;
        RECT 1.6500 0.4875 1.7100 0.5475 ;
        RECT 1.5450 0.1650 1.6050 0.2250 ;
        RECT 1.5450 0.7425 1.6050 0.8025 ;
        RECT 1.4400 0.4875 1.5000 0.5475 ;
        RECT 1.3350 0.2400 1.3950 0.3000 ;
        RECT 1.3350 0.8325 1.3950 0.8925 ;
        RECT 1.2300 0.4875 1.2900 0.5475 ;
        RECT 1.1250 0.3075 1.1850 0.3675 ;
        RECT 1.1250 0.7425 1.1850 0.8025 ;
        RECT 1.0200 0.4875 1.0800 0.5475 ;
        RECT 0.9150 0.1575 0.9750 0.2175 ;
        RECT 0.9150 0.8325 0.9750 0.8925 ;
        RECT 0.7050 0.1575 0.7650 0.2175 ;
        RECT 0.7050 0.8325 0.7650 0.8925 ;
        RECT 0.6000 0.4875 0.6600 0.5475 ;
        RECT 0.4950 0.2700 0.5550 0.3300 ;
        RECT 0.4950 0.7425 0.5550 0.8025 ;
        RECT 0.3900 0.4875 0.4500 0.5475 ;
        RECT 0.2850 0.1350 0.3450 0.1950 ;
        RECT 0.2850 0.8625 0.3450 0.9225 ;
        RECT 0.1800 0.4800 0.2400 0.5400 ;
        RECT 0.0750 0.2550 0.1350 0.3150 ;
        RECT 0.0750 0.7425 0.1350 0.8025 ;
        LAYER M1 ;
        RECT 2.3100 0.4500 2.3850 0.6825 ;
        RECT 2.0700 0.4500 2.3100 0.5700 ;
        RECT 1.6350 0.1500 2.2650 0.2250 ;
        RECT 1.7250 0.3000 1.8450 0.4050 ;
        RECT 1.5225 0.4800 1.7400 0.5700 ;
        RECT 1.4025 0.3150 1.7250 0.3900 ;
        RECT 1.5150 0.1500 1.6350 0.2400 ;
        RECT 1.4025 0.4650 1.5225 0.5700 ;
        RECT 1.3275 0.1500 1.4025 0.3900 ;
        RECT 0.8850 0.1500 1.3275 0.2250 ;
        RECT 0.9975 0.4650 1.3125 0.5700 ;
        RECT 0.9225 0.3000 1.2150 0.3750 ;
        RECT 0.8400 0.3000 0.9225 0.3975 ;
        RECT 0.5625 0.3225 0.8400 0.3975 ;
        RECT 0.4050 0.4800 0.6900 0.5550 ;
        RECT 0.4875 0.2400 0.5625 0.3975 ;
        RECT 0.3300 0.2700 0.4050 0.7875 ;
        RECT 0.1425 0.2700 0.3300 0.3450 ;
        RECT 0.1425 0.7125 0.3300 0.7875 ;
        RECT 0.0900 0.4200 0.2550 0.6375 ;
        RECT 0.0675 0.2250 0.1425 0.3450 ;
        RECT 0.0675 0.7125 0.1425 0.8325 ;
    END
END IND4_0011


MACRO IND4_0111
    CLASS CORE ;
    FOREIGN IND4_0111 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.2000 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 3.5175 0.2625 3.8325 0.7800 ;
        VIA 3.6750 0.3450 VIA12_slot ;
        VIA 3.6750 0.6975 VIA12_slot ;
        END
    END ZN
    PIN B3
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 3.2550 0.4125 3.3300 0.6075 ;
        RECT 2.7900 0.4125 3.2550 0.4875 ;
        VIA 3.2925 0.5250 VIA12_square ;
        END
    END B3
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 2.3775 0.4125 2.4525 0.6000 ;
        RECT 1.9125 0.4125 2.3775 0.4875 ;
        VIA 2.4150 0.5100 VIA12_square ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.5375 0.4125 1.6125 0.6000 ;
        RECT 1.0725 0.4125 1.5375 0.4875 ;
        VIA 1.5750 0.5100 VIA12_square ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.0900 0.5625 0.5550 0.6375 ;
        VIA 0.1725 0.6000 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.2000 -0.0750 4.2000 0.0750 ;
        RECT 1.0950 -0.0750 1.2000 0.2475 ;
        RECT 0.7875 -0.0750 1.0950 0.0750 ;
        RECT 0.6825 -0.0750 0.7875 0.2400 ;
        RECT 0.3750 -0.0750 0.6825 0.0750 ;
        RECT 0.2550 -0.0750 0.3750 0.1950 ;
        RECT 0.0000 -0.0750 0.2550 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 4.1325 0.9750 4.2000 1.1250 ;
        RECT 4.0575 0.7875 4.1325 1.1250 ;
        RECT 3.7350 0.9750 4.0575 1.1250 ;
        RECT 3.6150 0.8250 3.7350 1.1250 ;
        RECT 3.3150 0.9750 3.6150 1.1250 ;
        RECT 3.1950 0.8250 3.3150 1.1250 ;
        RECT 3.1050 0.9750 3.1950 1.1250 ;
        RECT 2.9850 0.8250 3.1050 1.1250 ;
        RECT 2.6850 0.9750 2.9850 1.1250 ;
        RECT 2.5650 0.8250 2.6850 1.1250 ;
        RECT 2.2650 0.9750 2.5650 1.1250 ;
        RECT 2.1450 0.8250 2.2650 1.1250 ;
        RECT 1.8450 0.9750 2.1450 1.1250 ;
        RECT 1.7250 0.8250 1.8450 1.1250 ;
        RECT 1.4250 0.9750 1.7250 1.1250 ;
        RECT 1.3050 0.8250 1.4250 1.1250 ;
        RECT 1.2150 0.9750 1.3050 1.1250 ;
        RECT 1.0950 0.8250 1.2150 1.1250 ;
        RECT 0.7950 0.9750 1.0950 1.1250 ;
        RECT 0.6750 0.8250 0.7950 1.1250 ;
        RECT 0.3750 0.9750 0.6750 1.1250 ;
        RECT 0.2550 0.8625 0.3750 1.1250 ;
        RECT 0.0000 0.9750 0.2550 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 4.0650 0.1725 4.1250 0.2325 ;
        RECT 4.0650 0.8175 4.1250 0.8775 ;
        RECT 3.9600 0.4950 4.0200 0.5550 ;
        RECT 3.8550 0.3225 3.9150 0.3825 ;
        RECT 3.8550 0.6675 3.9150 0.7275 ;
        RECT 3.7500 0.4950 3.8100 0.5550 ;
        RECT 3.6450 0.1575 3.7050 0.2175 ;
        RECT 3.6450 0.8325 3.7050 0.8925 ;
        RECT 3.5400 0.4950 3.6000 0.5550 ;
        RECT 3.4350 0.3225 3.4950 0.3825 ;
        RECT 3.4350 0.6675 3.4950 0.7275 ;
        RECT 3.3300 0.4950 3.3900 0.5550 ;
        RECT 3.2250 0.2325 3.2850 0.2925 ;
        RECT 3.2250 0.8325 3.2850 0.8925 ;
        RECT 3.0150 0.1575 3.0750 0.2175 ;
        RECT 3.0150 0.8325 3.0750 0.8925 ;
        RECT 2.9100 0.4800 2.9700 0.5400 ;
        RECT 2.8050 0.3075 2.8650 0.3675 ;
        RECT 2.8050 0.6675 2.8650 0.7275 ;
        RECT 2.7000 0.4800 2.7600 0.5400 ;
        RECT 2.5950 0.1575 2.6550 0.2175 ;
        RECT 2.5950 0.8325 2.6550 0.8925 ;
        RECT 2.4900 0.4800 2.5500 0.5400 ;
        RECT 2.3850 0.3075 2.4450 0.3675 ;
        RECT 2.3850 0.6675 2.4450 0.7275 ;
        RECT 2.2800 0.4800 2.3400 0.5400 ;
        RECT 2.1750 0.1575 2.2350 0.2175 ;
        RECT 2.1750 0.8325 2.2350 0.8925 ;
        RECT 2.0700 0.4800 2.1300 0.5400 ;
        RECT 1.9650 0.3075 2.0250 0.3675 ;
        RECT 1.9650 0.6675 2.0250 0.7275 ;
        RECT 1.8600 0.4800 1.9200 0.5400 ;
        RECT 1.7550 0.1575 1.8150 0.2175 ;
        RECT 1.7550 0.8325 1.8150 0.8925 ;
        RECT 1.6500 0.4800 1.7100 0.5400 ;
        RECT 1.5450 0.3075 1.6050 0.3675 ;
        RECT 1.5450 0.6675 1.6050 0.7275 ;
        RECT 1.4400 0.4800 1.5000 0.5400 ;
        RECT 1.3350 0.1575 1.3950 0.2175 ;
        RECT 1.3350 0.8325 1.3950 0.8925 ;
        RECT 1.1250 0.1575 1.1850 0.2175 ;
        RECT 1.1250 0.8325 1.1850 0.8925 ;
        RECT 1.0200 0.4950 1.0800 0.5550 ;
        RECT 0.9150 0.3225 0.9750 0.3825 ;
        RECT 0.9150 0.6675 0.9750 0.7275 ;
        RECT 0.8100 0.4950 0.8700 0.5550 ;
        RECT 0.7050 0.1575 0.7650 0.2175 ;
        RECT 0.7050 0.8325 0.7650 0.8925 ;
        RECT 0.6000 0.4950 0.6600 0.5550 ;
        RECT 0.4950 0.3075 0.5550 0.3675 ;
        RECT 0.4950 0.6900 0.5550 0.7500 ;
        RECT 0.3900 0.4950 0.4500 0.5550 ;
        RECT 0.2850 0.1350 0.3450 0.1950 ;
        RECT 0.2850 0.8625 0.3450 0.9225 ;
        RECT 0.1800 0.4800 0.2400 0.5400 ;
        RECT 0.0750 0.2550 0.1350 0.3150 ;
        RECT 0.0750 0.7425 0.1350 0.8025 ;
        LAYER M1 ;
        RECT 4.0425 0.1500 4.1475 0.2625 ;
        RECT 3.2100 0.4875 4.0650 0.5625 ;
        RECT 3.2925 0.1500 4.0425 0.2250 ;
        RECT 0.5625 0.6450 3.9450 0.7500 ;
        RECT 3.4125 0.3000 3.9375 0.4050 ;
        RECT 3.2175 0.1500 3.2925 0.3750 ;
        RECT 2.3550 0.3000 3.2175 0.3750 ;
        RECT 1.3050 0.1500 3.1050 0.2250 ;
        RECT 2.2575 0.4575 2.9925 0.5625 ;
        RECT 1.4175 0.4575 2.1525 0.5625 ;
        RECT 1.3425 0.3000 2.0550 0.3750 ;
        RECT 1.2600 0.3000 1.3425 0.3975 ;
        RECT 0.5625 0.3225 1.2600 0.3975 ;
        RECT 0.4050 0.4875 1.1100 0.5625 ;
        RECT 0.4875 0.2625 0.5625 0.3975 ;
        RECT 0.4875 0.6450 0.5625 0.8025 ;
        RECT 0.3300 0.2700 0.4050 0.7875 ;
        RECT 0.1425 0.2700 0.3300 0.3450 ;
        RECT 0.1425 0.7125 0.3300 0.7875 ;
        RECT 0.0900 0.4200 0.2550 0.6375 ;
        RECT 0.0675 0.2250 0.1425 0.3450 ;
        RECT 0.0675 0.7125 0.1425 0.8325 ;
    END
END IND4_0111


MACRO IND4_1000
    CLASS CORE ;
    FOREIGN IND4_1000 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.2600 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 1.1475 0.1500 1.2225 0.7425 ;
        RECT 1.1175 0.1500 1.1475 0.3825 ;
        RECT 0.9825 0.6675 1.1475 0.7425 ;
        RECT 0.9075 0.6675 0.9825 0.8700 ;
        RECT 0.5625 0.6675 0.9075 0.7425 ;
        RECT 0.4875 0.6675 0.5625 0.8700 ;
        END
    END ZN
    PIN B3
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.7275 0.2625 1.1925 0.3375 ;
        VIA 0.9975 0.3000 VIA12_square ;
        END
    END B3
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.4350 0.4125 0.9000 0.4875 ;
        VIA 0.7800 0.4500 VIA12_square ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.1425 0.2625 0.6075 0.3375 ;
        VIA 0.5250 0.3000 VIA12_square ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.0900 0.5625 0.5550 0.6375 ;
        VIA 0.1725 0.6000 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.3750 -0.0750 1.2600 0.0750 ;
        RECT 0.2550 -0.0750 0.3750 0.2025 ;
        RECT 0.0000 -0.0750 0.2550 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.2150 0.9750 1.2600 1.1250 ;
        RECT 1.0950 0.8325 1.2150 1.1250 ;
        RECT 0.7950 0.9750 1.0950 1.1250 ;
        RECT 0.6750 0.8400 0.7950 1.1250 ;
        RECT 0.3750 0.9750 0.6750 1.1250 ;
        RECT 0.2550 0.8625 0.3750 1.1250 ;
        RECT 0.0000 0.9750 0.2550 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.1250 0.1800 1.1850 0.2400 ;
        RECT 1.1250 0.8325 1.1850 0.8925 ;
        RECT 1.0125 0.4800 1.0725 0.5400 ;
        RECT 0.9150 0.7800 0.9750 0.8400 ;
        RECT 0.8100 0.4725 0.8700 0.5325 ;
        RECT 0.7050 0.8700 0.7650 0.9300 ;
        RECT 0.6000 0.4650 0.6600 0.5250 ;
        RECT 0.4950 0.7800 0.5550 0.8400 ;
        RECT 0.3900 0.4800 0.4500 0.5400 ;
        RECT 0.2850 0.1275 0.3450 0.1875 ;
        RECT 0.2850 0.8700 0.3450 0.9300 ;
        RECT 0.1800 0.4800 0.2400 0.5400 ;
        RECT 0.0750 0.1725 0.1350 0.2325 ;
        RECT 0.0750 0.8175 0.1350 0.8775 ;
        LAYER M1 ;
        RECT 1.0425 0.4500 1.0725 0.5700 ;
        RECT 0.9600 0.2175 1.0425 0.5700 ;
        RECT 0.8325 0.4425 0.8700 0.5925 ;
        RECT 0.7425 0.2775 0.8325 0.5925 ;
        RECT 0.5775 0.2175 0.6675 0.5625 ;
        RECT 0.4875 0.2175 0.5775 0.3825 ;
        RECT 0.4125 0.4575 0.4725 0.5625 ;
        RECT 0.3375 0.2775 0.4125 0.7875 ;
        RECT 0.1575 0.2775 0.3375 0.3525 ;
        RECT 0.1575 0.7125 0.3375 0.7875 ;
        RECT 0.0900 0.4275 0.2550 0.6375 ;
        RECT 0.0525 0.1500 0.1575 0.3525 ;
        RECT 0.0525 0.7125 0.1575 0.9000 ;
    END
END IND4_1000


MACRO IND4_1010
    CLASS CORE ;
    FOREIGN IND4_1010 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.2600 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 1.1475 0.2175 1.2225 0.7425 ;
        RECT 1.1175 0.2175 1.1475 0.3825 ;
        RECT 0.5625 0.6675 1.1475 0.7425 ;
        RECT 0.4875 0.6675 0.5625 0.8325 ;
        END
    END ZN
    PIN B3
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.7275 0.2625 1.1925 0.3375 ;
        VIA 0.9975 0.3000 VIA12_square ;
        END
    END B3
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.4350 0.4125 0.9000 0.4875 ;
        VIA 0.7800 0.4500 VIA12_square ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.1425 0.2625 0.6075 0.3375 ;
        VIA 0.5250 0.3000 VIA12_square ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.0900 0.5625 0.5550 0.6375 ;
        VIA 0.1725 0.6000 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.3750 -0.0750 1.2600 0.0750 ;
        RECT 0.2550 -0.0750 0.3750 0.2025 ;
        RECT 0.0000 -0.0750 0.2550 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.2150 0.9750 1.2600 1.1250 ;
        RECT 1.0950 0.8325 1.2150 1.1250 ;
        RECT 0.7950 0.9750 1.0950 1.1250 ;
        RECT 0.6750 0.8400 0.7950 1.1250 ;
        RECT 0.3750 0.9750 0.6750 1.1250 ;
        RECT 0.2550 0.8625 0.3750 1.1250 ;
        RECT 0.0000 0.9750 0.2550 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.1250 0.2700 1.1850 0.3300 ;
        RECT 1.1250 0.8325 1.1850 0.8925 ;
        RECT 1.0125 0.4800 1.0725 0.5400 ;
        RECT 0.9150 0.6750 0.9750 0.7350 ;
        RECT 0.8100 0.4725 0.8700 0.5325 ;
        RECT 0.7050 0.8700 0.7650 0.9300 ;
        RECT 0.6000 0.4650 0.6600 0.5250 ;
        RECT 0.4950 0.7275 0.5550 0.7875 ;
        RECT 0.3900 0.4800 0.4500 0.5400 ;
        RECT 0.2850 0.1275 0.3450 0.1875 ;
        RECT 0.2850 0.8700 0.3450 0.9300 ;
        RECT 0.1800 0.4800 0.2400 0.5400 ;
        RECT 0.0750 0.2250 0.1350 0.2850 ;
        RECT 0.0750 0.7500 0.1350 0.8100 ;
        LAYER M1 ;
        RECT 1.0425 0.4500 1.0725 0.5700 ;
        RECT 0.9600 0.2175 1.0425 0.5700 ;
        RECT 0.8325 0.4425 0.8700 0.5925 ;
        RECT 0.7425 0.2775 0.8325 0.5925 ;
        RECT 0.5775 0.2175 0.6675 0.5625 ;
        RECT 0.4875 0.2175 0.5775 0.3825 ;
        RECT 0.4125 0.4575 0.4725 0.5625 ;
        RECT 0.3375 0.2775 0.4125 0.7875 ;
        RECT 0.1425 0.2775 0.3375 0.3525 ;
        RECT 0.1425 0.7125 0.3375 0.7875 ;
        RECT 0.0900 0.4275 0.2550 0.6375 ;
        RECT 0.0675 0.1800 0.1425 0.3525 ;
        RECT 0.0675 0.7125 0.1425 0.8400 ;
    END
END IND4_1010


MACRO INR2_0010
    CLASS CORE ;
    FOREIGN INR2_0010 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.2500 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 2.3625 0.2850 2.5200 0.4050 ;
        RECT 2.3625 0.6375 2.5200 0.7575 ;
        RECT 2.0475 0.2850 2.3625 0.7575 ;
        RECT 1.8900 0.2850 2.0475 0.4050 ;
        RECT 1.8900 0.6375 2.0475 0.7575 ;
        VIA 2.3625 0.3450 VIA12_slot ;
        VIA 2.3625 0.6975 VIA12_slot ;
        VIA 2.0475 0.3450 VIA12_slot ;
        VIA 2.0475 0.6975 VIA12_slot ;
        END
    END ZN
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 4.9125 0.4125 5.0775 0.6375 ;
        RECT 2.6700 0.4950 4.9125 0.6375 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1425 0.4500 0.6600 0.5700 ;
        RECT 0.0675 0.3675 0.1425 0.6825 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 5.1825 -0.0750 5.2500 0.0750 ;
        RECT 5.1075 -0.0750 5.1825 0.2700 ;
        RECT 4.7850 -0.0750 5.1075 0.0750 ;
        RECT 4.6650 -0.0750 4.7850 0.1875 ;
        RECT 4.3650 -0.0750 4.6650 0.0750 ;
        RECT 4.2450 -0.0750 4.3650 0.1875 ;
        RECT 3.9450 -0.0750 4.2450 0.0750 ;
        RECT 3.8250 -0.0750 3.9450 0.1875 ;
        RECT 3.5250 -0.0750 3.8250 0.0750 ;
        RECT 3.4050 -0.0750 3.5250 0.1875 ;
        RECT 3.1050 -0.0750 3.4050 0.0750 ;
        RECT 2.9850 -0.0750 3.1050 0.1875 ;
        RECT 2.6850 -0.0750 2.9850 0.0750 ;
        RECT 2.5650 -0.0750 2.6850 0.1875 ;
        RECT 2.2650 -0.0750 2.5650 0.0750 ;
        RECT 2.1450 -0.0750 2.2650 0.1875 ;
        RECT 1.8450 -0.0750 2.1450 0.0750 ;
        RECT 1.7250 -0.0750 1.8450 0.1875 ;
        RECT 1.4250 -0.0750 1.7250 0.0750 ;
        RECT 1.3050 -0.0750 1.4250 0.1875 ;
        RECT 0.9975 -0.0750 1.3050 0.0750 ;
        RECT 0.8925 -0.0750 0.9975 0.2625 ;
        RECT 0.5850 -0.0750 0.8925 0.0750 ;
        RECT 0.4650 -0.0750 0.5850 0.1950 ;
        RECT 0.1575 -0.0750 0.4650 0.0750 ;
        RECT 0.0525 -0.0750 0.1575 0.2625 ;
        RECT 0.0000 -0.0750 0.0525 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 4.9950 0.9750 5.2500 1.1250 ;
        RECT 4.8750 0.8625 4.9950 1.1250 ;
        RECT 4.5750 0.9750 4.8750 1.1250 ;
        RECT 4.4550 0.8625 4.5750 1.1250 ;
        RECT 4.1550 0.9750 4.4550 1.1250 ;
        RECT 4.0350 0.8625 4.1550 1.1250 ;
        RECT 3.7350 0.9750 4.0350 1.1250 ;
        RECT 3.6150 0.8625 3.7350 1.1250 ;
        RECT 3.3150 0.9750 3.6150 1.1250 ;
        RECT 3.1950 0.8625 3.3150 1.1250 ;
        RECT 2.8950 0.9750 3.1950 1.1250 ;
        RECT 2.7750 0.8625 2.8950 1.1250 ;
        RECT 0.5850 0.9750 2.7750 1.1250 ;
        RECT 0.4650 0.8250 0.5850 1.1250 ;
        RECT 0.1575 0.9750 0.4650 1.1250 ;
        RECT 0.0525 0.7875 0.1575 1.1250 ;
        RECT 0.0000 0.9750 0.0525 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 5.1150 0.1575 5.1750 0.2175 ;
        RECT 5.1150 0.7800 5.1750 0.8400 ;
        RECT 5.0100 0.4950 5.0700 0.5550 ;
        RECT 4.9050 0.1725 4.9650 0.2325 ;
        RECT 4.9050 0.8625 4.9650 0.9225 ;
        RECT 4.8000 0.4950 4.8600 0.5550 ;
        RECT 4.6950 0.1275 4.7550 0.1875 ;
        RECT 4.6950 0.7200 4.7550 0.7800 ;
        RECT 4.5900 0.4950 4.6500 0.5550 ;
        RECT 4.4850 0.1725 4.5450 0.2325 ;
        RECT 4.4850 0.8625 4.5450 0.9225 ;
        RECT 4.3800 0.4950 4.4400 0.5550 ;
        RECT 4.2750 0.1275 4.3350 0.1875 ;
        RECT 4.2750 0.7200 4.3350 0.7800 ;
        RECT 4.1700 0.4950 4.2300 0.5550 ;
        RECT 4.0650 0.1725 4.1250 0.2325 ;
        RECT 4.0650 0.8625 4.1250 0.9225 ;
        RECT 3.9600 0.4950 4.0200 0.5550 ;
        RECT 3.8550 0.1275 3.9150 0.1875 ;
        RECT 3.8550 0.7200 3.9150 0.7800 ;
        RECT 3.7500 0.4950 3.8100 0.5550 ;
        RECT 3.6450 0.1725 3.7050 0.2325 ;
        RECT 3.6450 0.8625 3.7050 0.9225 ;
        RECT 3.5400 0.4950 3.6000 0.5550 ;
        RECT 3.4350 0.1275 3.4950 0.1875 ;
        RECT 3.4350 0.7200 3.4950 0.7800 ;
        RECT 3.3300 0.4950 3.3900 0.5550 ;
        RECT 3.2250 0.2925 3.2850 0.3525 ;
        RECT 3.2250 0.8625 3.2850 0.9225 ;
        RECT 3.1200 0.4950 3.1800 0.5550 ;
        RECT 3.0150 0.1275 3.0750 0.1875 ;
        RECT 3.0150 0.7200 3.0750 0.7800 ;
        RECT 2.9100 0.4950 2.9700 0.5550 ;
        RECT 2.8050 0.2925 2.8650 0.3525 ;
        RECT 2.8050 0.8625 2.8650 0.9225 ;
        RECT 2.7000 0.4950 2.7600 0.5550 ;
        RECT 2.5950 0.1275 2.6550 0.1875 ;
        RECT 2.5950 0.8325 2.6550 0.8925 ;
        RECT 2.4900 0.4800 2.5500 0.5400 ;
        RECT 2.3850 0.2925 2.4450 0.3525 ;
        RECT 2.3850 0.6900 2.4450 0.7500 ;
        RECT 2.2800 0.4800 2.3400 0.5400 ;
        RECT 2.1750 0.1275 2.2350 0.1875 ;
        RECT 2.1750 0.8325 2.2350 0.8925 ;
        RECT 2.0700 0.4800 2.1300 0.5400 ;
        RECT 1.9650 0.2925 2.0250 0.3525 ;
        RECT 1.9650 0.6900 2.0250 0.7500 ;
        RECT 1.8600 0.4800 1.9200 0.5400 ;
        RECT 1.7550 0.1275 1.8150 0.1875 ;
        RECT 1.7550 0.8325 1.8150 0.8925 ;
        RECT 1.6500 0.4800 1.7100 0.5400 ;
        RECT 1.5450 0.2925 1.6050 0.3525 ;
        RECT 1.5450 0.6900 1.6050 0.7500 ;
        RECT 1.4400 0.4800 1.5000 0.5400 ;
        RECT 1.3350 0.1275 1.3950 0.1875 ;
        RECT 1.3350 0.8325 1.3950 0.8925 ;
        RECT 1.2300 0.4800 1.2900 0.5400 ;
        RECT 1.1250 0.2925 1.1850 0.3525 ;
        RECT 1.1250 0.6900 1.1850 0.7500 ;
        RECT 1.0200 0.4800 1.0800 0.5400 ;
        RECT 0.9150 0.1725 0.9750 0.2325 ;
        RECT 0.9150 0.8100 0.9750 0.8700 ;
        RECT 0.7050 0.2925 0.7650 0.3525 ;
        RECT 0.7050 0.6900 0.7650 0.7500 ;
        RECT 0.6000 0.4800 0.6600 0.5400 ;
        RECT 0.4950 0.1275 0.5550 0.1875 ;
        RECT 0.4950 0.8250 0.5550 0.8850 ;
        RECT 0.3900 0.4800 0.4500 0.5400 ;
        RECT 0.2850 0.2925 0.3450 0.3525 ;
        RECT 0.2850 0.6975 0.3450 0.7575 ;
        RECT 0.1800 0.4800 0.2400 0.5400 ;
        RECT 0.0750 0.1725 0.1350 0.2325 ;
        RECT 0.0750 0.8175 0.1350 0.8775 ;
        LAYER M1 ;
        RECT 5.1075 0.7125 5.1825 0.8700 ;
        RECT 2.6925 0.7125 5.1075 0.7875 ;
        RECT 4.8825 0.1500 4.9875 0.3375 ;
        RECT 4.8375 0.2625 4.8825 0.3375 ;
        RECT 4.5675 0.2625 4.8375 0.3825 ;
        RECT 4.4625 0.1500 4.5675 0.3825 ;
        RECT 4.1475 0.2625 4.4625 0.3825 ;
        RECT 4.0425 0.1500 4.1475 0.3825 ;
        RECT 3.7275 0.2625 4.0425 0.3825 ;
        RECT 3.6225 0.1500 3.7275 0.3825 ;
        RECT 1.1175 0.2625 3.6225 0.3825 ;
        RECT 2.6175 0.7125 2.6925 0.9000 ;
        RECT 0.9975 0.8250 2.6175 0.9000 ;
        RECT 0.8100 0.4650 2.5800 0.5700 ;
        RECT 1.0950 0.6450 2.5425 0.7500 ;
        RECT 0.8925 0.7800 0.9975 0.9000 ;
        RECT 0.7350 0.2700 0.8100 0.7500 ;
        RECT 0.2550 0.2700 0.7350 0.3750 ;
        RECT 0.3750 0.6750 0.7350 0.7500 ;
        RECT 0.2625 0.6750 0.3750 0.7800 ;
        LAYER M2 ;
        RECT 2.3925 0.2850 2.5200 0.4050 ;
        RECT 2.3925 0.6375 2.5200 0.7575 ;
        RECT 1.8900 0.2850 2.0175 0.4050 ;
        RECT 1.8900 0.6375 2.0175 0.7575 ;
    END
END INR2_0010


MACRO INR2_0011
    CLASS CORE ;
    FOREIGN INR2_0011 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.2600 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 0.9075 0.1125 0.9975 0.1875 ;
        RECT 0.8325 0.1125 0.9075 0.9375 ;
        RECT 0.3675 0.8625 0.8325 0.9375 ;
        VIA 0.8700 0.3450 VIA12_square ;
        VIA 0.8700 0.8475 VIA12_square ;
        END
    END ZN
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.6825 0.1125 0.7575 0.6900 ;
        RECT 0.2175 0.1125 0.6825 0.1875 ;
        VIA 0.7200 0.5100 VIA12_square ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.0975 0.5625 0.5625 0.6375 ;
        VIA 0.1800 0.6000 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.2000 -0.0750 1.2600 0.0750 ;
        RECT 1.1250 -0.0750 1.2000 0.2475 ;
        RECT 0.7875 -0.0750 1.1250 0.0750 ;
        RECT 0.6825 -0.0750 0.7875 0.2250 ;
        RECT 0.3750 -0.0750 0.6825 0.0750 ;
        RECT 0.2550 -0.0750 0.3750 0.1875 ;
        RECT 0.0000 -0.0750 0.2550 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.2075 0.9750 1.2600 1.1250 ;
        RECT 1.1025 0.8100 1.2075 1.1250 ;
        RECT 0.3750 0.9750 1.1025 1.1250 ;
        RECT 0.2550 0.8625 0.3750 1.1250 ;
        RECT 0.0000 0.9750 0.2550 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.1250 0.1575 1.1850 0.2175 ;
        RECT 1.1250 0.8325 1.1850 0.8925 ;
        RECT 1.0200 0.4950 1.0800 0.5550 ;
        RECT 0.9150 0.2475 0.9750 0.3075 ;
        RECT 0.8100 0.4950 0.8700 0.5550 ;
        RECT 0.7050 0.1425 0.7650 0.2025 ;
        RECT 0.7050 0.8175 0.7650 0.8775 ;
        RECT 0.6000 0.4950 0.6600 0.5550 ;
        RECT 0.4950 0.2475 0.5550 0.3075 ;
        RECT 0.3900 0.4800 0.4500 0.5400 ;
        RECT 0.2850 0.1275 0.3450 0.1875 ;
        RECT 0.2850 0.8625 0.3450 0.9225 ;
        RECT 0.1800 0.4800 0.2400 0.5400 ;
        RECT 0.0750 0.2475 0.1350 0.3075 ;
        RECT 0.0750 0.7425 0.1350 0.8025 ;
        LAYER M1 ;
        RECT 1.0425 0.4725 1.1025 0.5775 ;
        RECT 0.9675 0.4725 1.0425 0.7275 ;
        RECT 0.6525 0.8025 0.9975 0.9000 ;
        RECT 0.9075 0.2025 0.9825 0.3825 ;
        RECT 0.4500 0.6525 0.9675 0.7275 ;
        RECT 0.5625 0.3075 0.9075 0.3825 ;
        RECT 0.5775 0.4725 0.8925 0.5775 ;
        RECT 0.4875 0.2025 0.5625 0.3825 ;
        RECT 0.4125 0.4500 0.4500 0.7275 ;
        RECT 0.3375 0.2625 0.4125 0.7875 ;
        RECT 0.1425 0.2625 0.3375 0.3375 ;
        RECT 0.1425 0.7125 0.3375 0.7875 ;
        RECT 0.0975 0.4125 0.2625 0.6375 ;
        RECT 0.0675 0.2175 0.1425 0.3375 ;
        RECT 0.0675 0.7125 0.1425 0.8325 ;
    END
END INR2_0011


MACRO INR2_0111
    CLASS CORE ;
    FOREIGN INR2_0111 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.1000 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 1.2075 0.2625 1.5225 0.7875 ;
        VIA 1.3650 0.3450 VIA12_slot ;
        VIA 1.3650 0.7050 VIA12_slot ;
        END
    END ZN
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.9825 0.2625 1.0575 0.6075 ;
        RECT 0.5625 0.2625 0.9825 0.3375 ;
        VIA 1.0200 0.5175 VIA12_square ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.0975 0.5625 0.5625 0.6375 ;
        VIA 0.1800 0.6000 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 2.0475 -0.0750 2.1000 0.0750 ;
        RECT 1.9425 -0.0750 2.0475 0.2700 ;
        RECT 1.6275 -0.0750 1.9425 0.0750 ;
        RECT 1.5225 -0.0750 1.6275 0.2100 ;
        RECT 1.2075 -0.0750 1.5225 0.0750 ;
        RECT 1.1025 -0.0750 1.2075 0.2100 ;
        RECT 0.7875 -0.0750 1.1025 0.0750 ;
        RECT 0.6825 -0.0750 0.7875 0.2100 ;
        RECT 0.3750 -0.0750 0.6825 0.0750 ;
        RECT 0.2550 -0.0750 0.3750 0.1950 ;
        RECT 0.0000 -0.0750 0.2550 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 2.0325 0.9750 2.1000 1.1250 ;
        RECT 1.9575 0.7875 2.0325 1.1250 ;
        RECT 0.7950 0.9750 1.9575 1.1250 ;
        RECT 0.6750 0.8400 0.7950 1.1250 ;
        RECT 0.3750 0.9750 0.6750 1.1250 ;
        RECT 0.2550 0.8700 0.3750 1.1250 ;
        RECT 0.0000 0.9750 0.2550 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.9650 0.1725 2.0250 0.2325 ;
        RECT 1.9650 0.8325 2.0250 0.8925 ;
        RECT 1.8600 0.4950 1.9200 0.5550 ;
        RECT 1.7550 0.3075 1.8150 0.3675 ;
        RECT 1.7550 0.8325 1.8150 0.8925 ;
        RECT 1.6500 0.4875 1.7100 0.5475 ;
        RECT 1.5450 0.1275 1.6050 0.1875 ;
        RECT 1.5450 0.6900 1.6050 0.7500 ;
        RECT 1.4400 0.4875 1.5000 0.5475 ;
        RECT 1.3350 0.3150 1.3950 0.3750 ;
        RECT 1.3350 0.8325 1.3950 0.8925 ;
        RECT 1.2300 0.4875 1.2900 0.5475 ;
        RECT 1.1250 0.1275 1.1850 0.1875 ;
        RECT 1.1250 0.6900 1.1850 0.7500 ;
        RECT 1.0200 0.4875 1.0800 0.5475 ;
        RECT 0.9150 0.3150 0.9750 0.3750 ;
        RECT 0.9150 0.7350 0.9750 0.7950 ;
        RECT 0.8025 0.4950 0.8625 0.5550 ;
        RECT 0.7050 0.1275 0.7650 0.1875 ;
        RECT 0.7050 0.8550 0.7650 0.9150 ;
        RECT 0.6000 0.4950 0.6600 0.5550 ;
        RECT 0.4950 0.2325 0.5550 0.2925 ;
        RECT 0.4950 0.7200 0.5550 0.7800 ;
        RECT 0.3900 0.4950 0.4500 0.5550 ;
        RECT 0.2850 0.1275 0.3450 0.1875 ;
        RECT 0.2850 0.8700 0.3450 0.9300 ;
        RECT 0.1800 0.4800 0.2400 0.5400 ;
        RECT 0.0750 0.2550 0.1350 0.3150 ;
        RECT 0.0750 0.7500 0.1350 0.8100 ;
        LAYER M1 ;
        RECT 1.8450 0.4650 2.0400 0.6375 ;
        RECT 0.9825 0.8250 1.8450 0.9000 ;
        RECT 1.7325 0.2850 1.8375 0.3900 ;
        RECT 1.0275 0.4800 1.7400 0.5550 ;
        RECT 0.9450 0.2850 1.7325 0.4050 ;
        RECT 1.0950 0.6600 1.7325 0.7500 ;
        RECT 0.9375 0.4800 1.0275 0.5850 ;
        RECT 0.9075 0.6900 0.9825 0.9000 ;
        RECT 0.5625 0.2850 0.9450 0.3900 ;
        RECT 0.5625 0.6900 0.9075 0.7650 ;
        RECT 0.4125 0.4650 0.8625 0.5850 ;
        RECT 0.4875 0.1950 0.5625 0.3900 ;
        RECT 0.4875 0.6900 0.5625 0.8100 ;
        RECT 0.3375 0.2700 0.4125 0.7950 ;
        RECT 0.1425 0.2700 0.3375 0.3450 ;
        RECT 0.1425 0.7200 0.3375 0.7950 ;
        RECT 0.0975 0.4200 0.2625 0.6450 ;
        RECT 0.0675 0.2250 0.1425 0.3450 ;
        RECT 0.0675 0.7200 0.1425 0.8400 ;
        LAYER VIA1 ;
        RECT 1.8900 0.5625 1.9650 0.6375 ;
        RECT 0.7125 0.4875 0.7875 0.5625 ;
        LAYER M2 ;
        RECT 1.7475 0.5625 2.0100 0.6375 ;
        RECT 1.6725 0.5625 1.7475 0.9375 ;
        RECT 0.7725 0.8625 1.6725 0.9375 ;
        RECT 0.7725 0.4425 0.8025 0.6075 ;
        RECT 0.6975 0.4425 0.7725 0.9375 ;
    END
END INR2_0111


MACRO INR2_1000
    CLASS CORE ;
    FOREIGN INR2_1000 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.8400 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.7275 0.3075 0.8025 0.9000 ;
        RECT 0.5625 0.3075 0.7275 0.3825 ;
        RECT 0.6750 0.8025 0.7275 0.9000 ;
        RECT 0.4875 0.1800 0.5625 0.3825 ;
        END
    END ZN
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.5625 0.4575 0.6525 0.7125 ;
        RECT 0.5475 0.4575 0.5625 0.8325 ;
        RECT 0.4875 0.6375 0.5475 0.8325 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.0975 0.4125 0.5625 0.4875 ;
        VIA 0.1800 0.4500 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.7950 -0.0750 0.8400 0.0750 ;
        RECT 0.6750 -0.0750 0.7950 0.2325 ;
        RECT 0.3750 -0.0750 0.6750 0.0750 ;
        RECT 0.2550 -0.0750 0.3750 0.1875 ;
        RECT 0.0000 -0.0750 0.2550 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.3750 0.9750 0.8400 1.1250 ;
        RECT 0.2550 0.8325 0.3750 1.1250 ;
        RECT 0.0000 0.9750 0.2550 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 0.7050 0.1575 0.7650 0.2175 ;
        RECT 0.7050 0.8175 0.7650 0.8775 ;
        RECT 0.5925 0.4950 0.6525 0.5550 ;
        RECT 0.4950 0.2100 0.5550 0.2700 ;
        RECT 0.3825 0.4875 0.4425 0.5475 ;
        RECT 0.2850 0.1200 0.3450 0.1800 ;
        RECT 0.2850 0.8400 0.3450 0.9000 ;
        RECT 0.1800 0.4875 0.2400 0.5475 ;
        RECT 0.0750 0.1725 0.1350 0.2325 ;
        RECT 0.0750 0.8175 0.1350 0.8775 ;
        LAYER M1 ;
        RECT 0.4125 0.4575 0.4425 0.5775 ;
        RECT 0.3375 0.2625 0.4125 0.7575 ;
        RECT 0.1575 0.2625 0.3375 0.3375 ;
        RECT 0.1575 0.6825 0.3375 0.7575 ;
        RECT 0.0975 0.4125 0.2625 0.6075 ;
        RECT 0.0525 0.1500 0.1575 0.3375 ;
        RECT 0.0525 0.6825 0.1575 0.9000 ;
    END
END INR2_1000


MACRO INR2_1010
    CLASS CORE ;
    FOREIGN INR2_1010 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.8400 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.7275 0.3075 0.8025 0.8850 ;
        RECT 0.5625 0.3075 0.7275 0.3825 ;
        RECT 0.6975 0.7650 0.7275 0.8850 ;
        RECT 0.4875 0.2175 0.5625 0.3825 ;
        END
    END ZN
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.6225 0.4575 0.6525 0.5925 ;
        RECT 0.5475 0.4575 0.6225 0.8325 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.2925 0.2625 0.3825 0.3900 ;
        RECT 0.2100 0.2625 0.2925 0.6075 ;
        RECT 0.1875 0.4500 0.2100 0.6075 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.7950 -0.0750 0.8400 0.0750 ;
        RECT 0.6750 -0.0750 0.7950 0.2325 ;
        RECT 0.3750 -0.0750 0.6750 0.0750 ;
        RECT 0.2550 -0.0750 0.3750 0.1875 ;
        RECT 0.0000 -0.0750 0.2550 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.3750 0.9750 0.8400 1.1250 ;
        RECT 0.2550 0.8325 0.3750 1.1250 ;
        RECT 0.0000 0.9750 0.2550 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 0.7050 0.1575 0.7650 0.2175 ;
        RECT 0.7050 0.7950 0.7650 0.8550 ;
        RECT 0.5925 0.4950 0.6525 0.5550 ;
        RECT 0.4950 0.2475 0.5550 0.3075 ;
        RECT 0.3900 0.4875 0.4500 0.5475 ;
        RECT 0.2850 0.1200 0.3450 0.1800 ;
        RECT 0.2850 0.8400 0.3450 0.9000 ;
        RECT 0.1875 0.4875 0.2475 0.5475 ;
        RECT 0.0750 0.2100 0.1350 0.2700 ;
        RECT 0.0750 0.6900 0.1350 0.7500 ;
        LAYER M1 ;
        RECT 0.4425 0.4650 0.4725 0.5700 ;
        RECT 0.3675 0.4650 0.4425 0.7575 ;
        RECT 0.1125 0.6825 0.3675 0.7575 ;
        RECT 0.1125 0.1800 0.1350 0.3000 ;
        RECT 0.0375 0.1800 0.1125 0.7575 ;
    END
END INR2_1010


MACRO INR3_0011
    CLASS CORE ;
    FOREIGN INR3_0011 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.8900 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 0.6900 0.2625 1.2450 0.3375 ;
        VIA 1.1550 0.3000 VIA12_square ;
        END
    END ZN
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.1025 0.4425 1.2075 0.6375 ;
        RECT 0.6525 0.5625 1.1025 0.6375 ;
        VIA 1.1550 0.5250 VIA12_square ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.7475 0.3675 1.8225 0.6825 ;
        RECT 1.3875 0.4650 1.7475 0.5700 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.0900 0.4125 0.5550 0.4875 ;
        VIA 0.1725 0.4500 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.8375 -0.0750 1.8900 0.0750 ;
        RECT 1.7325 -0.0750 1.8375 0.2400 ;
        RECT 1.4250 -0.0750 1.7325 0.0750 ;
        RECT 1.3050 -0.0750 1.4250 0.2250 ;
        RECT 1.0050 -0.0750 1.3050 0.0750 ;
        RECT 0.8850 -0.0750 1.0050 0.2250 ;
        RECT 0.7950 -0.0750 0.8850 0.0750 ;
        RECT 0.6750 -0.0750 0.7950 0.2250 ;
        RECT 0.3750 -0.0750 0.6750 0.0750 ;
        RECT 0.2550 -0.0750 0.3750 0.1875 ;
        RECT 0.0000 -0.0750 0.2550 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.7800 0.9750 1.8900 1.1250 ;
        RECT 0.6750 0.8025 0.7800 1.1250 ;
        RECT 0.3750 0.9750 0.6750 1.1250 ;
        RECT 0.2550 0.8550 0.3750 1.1250 ;
        RECT 0.0000 0.9750 0.2550 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.7550 0.1575 1.8150 0.2175 ;
        RECT 1.7550 0.8175 1.8150 0.8775 ;
        RECT 1.6500 0.4800 1.7100 0.5400 ;
        RECT 1.5450 0.2775 1.6050 0.3375 ;
        RECT 1.5450 0.6750 1.6050 0.7350 ;
        RECT 1.4400 0.4800 1.5000 0.5400 ;
        RECT 1.3350 0.1575 1.3950 0.2175 ;
        RECT 1.3350 0.8325 1.3950 0.8925 ;
        RECT 1.2300 0.4950 1.2900 0.5550 ;
        RECT 1.1250 0.2775 1.1850 0.3375 ;
        RECT 1.1250 0.6825 1.1850 0.7425 ;
        RECT 1.0200 0.4950 1.0800 0.5550 ;
        RECT 0.9150 0.1575 0.9750 0.2175 ;
        RECT 0.9150 0.8325 0.9750 0.8925 ;
        RECT 0.7050 0.1575 0.7650 0.2175 ;
        RECT 0.7050 0.8325 0.7650 0.8925 ;
        RECT 0.6000 0.4950 0.6600 0.5550 ;
        RECT 0.4950 0.2775 0.5550 0.3375 ;
        RECT 0.4950 0.6975 0.5550 0.7575 ;
        RECT 0.3900 0.4950 0.4500 0.5550 ;
        RECT 0.2850 0.1200 0.3450 0.1800 ;
        RECT 0.2850 0.8550 0.3450 0.9150 ;
        RECT 0.1800 0.4800 0.2400 0.5400 ;
        RECT 0.0750 0.2475 0.1350 0.3075 ;
        RECT 0.0750 0.7350 0.1350 0.7950 ;
        LAYER M1 ;
        RECT 1.7325 0.7950 1.8375 0.9000 ;
        RECT 0.8850 0.8250 1.7325 0.9000 ;
        RECT 1.4250 0.6450 1.6725 0.7500 ;
        RECT 1.5375 0.2175 1.6125 0.3900 ;
        RECT 1.1925 0.3150 1.5375 0.3900 ;
        RECT 1.3200 0.6600 1.4250 0.7500 ;
        RECT 0.9975 0.4725 1.3125 0.5775 ;
        RECT 0.9225 0.6750 1.2150 0.7500 ;
        RECT 1.1175 0.2175 1.1925 0.3900 ;
        RECT 0.9225 0.3150 1.1175 0.3900 ;
        RECT 0.8400 0.3150 0.9225 0.7500 ;
        RECT 0.5625 0.3150 0.8400 0.3900 ;
        RECT 0.6000 0.6525 0.7350 0.7275 ;
        RECT 0.4050 0.4875 0.6900 0.5625 ;
        RECT 0.4875 0.6525 0.6000 0.9000 ;
        RECT 0.4875 0.2175 0.5625 0.3900 ;
        RECT 0.3300 0.2625 0.4050 0.7800 ;
        RECT 0.1425 0.2625 0.3300 0.3375 ;
        RECT 0.1425 0.7050 0.3300 0.7800 ;
        RECT 0.0900 0.4125 0.2550 0.6300 ;
        RECT 0.0675 0.2175 0.1425 0.3375 ;
        RECT 0.0675 0.7050 0.1425 0.8250 ;
        LAYER VIA1 ;
        RECT 1.3725 0.6750 1.4475 0.7500 ;
        RECT 0.5100 0.7125 0.5850 0.7875 ;
        LAYER M2 ;
        RECT 1.3800 0.6750 1.4925 0.7500 ;
        RECT 1.3050 0.6750 1.3800 0.7875 ;
        RECT 0.4425 0.7125 1.3050 0.7875 ;
    END
END INR3_0011


MACRO INR3_0111
    CLASS CORE ;
    FOREIGN INR3_0111 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.1500 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 2.4675 0.2625 2.7825 0.7800 ;
        VIA 2.6250 0.3450 VIA12_slot ;
        VIA 2.6250 0.6975 VIA12_slot ;
        END
    END ZN
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 3.0075 0.3675 3.0825 0.6825 ;
        RECT 2.2575 0.4725 3.0075 0.5775 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.7475 0.4125 1.8225 0.6075 ;
        RECT 1.2825 0.4125 1.7475 0.4875 ;
        VIA 1.7850 0.5250 VIA12_square ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.0900 0.4125 0.5550 0.4875 ;
        VIA 0.1725 0.4500 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 3.0825 -0.0750 3.1500 0.0750 ;
        RECT 3.0075 -0.0750 3.0825 0.2625 ;
        RECT 2.6850 -0.0750 3.0075 0.0750 ;
        RECT 2.5650 -0.0750 2.6850 0.2175 ;
        RECT 2.2650 -0.0750 2.5650 0.0750 ;
        RECT 2.1450 -0.0750 2.2650 0.2175 ;
        RECT 1.8450 -0.0750 2.1450 0.0750 ;
        RECT 1.7250 -0.0750 1.8450 0.2175 ;
        RECT 1.4250 -0.0750 1.7250 0.0750 ;
        RECT 1.3050 -0.0750 1.4250 0.2175 ;
        RECT 1.2150 -0.0750 1.3050 0.0750 ;
        RECT 1.0950 -0.0750 1.2150 0.2175 ;
        RECT 0.7950 -0.0750 1.0950 0.0750 ;
        RECT 0.6750 -0.0750 0.7950 0.2175 ;
        RECT 0.3750 -0.0750 0.6750 0.0750 ;
        RECT 0.2550 -0.0750 0.3750 0.1875 ;
        RECT 0.0000 -0.0750 0.2550 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.2000 0.9750 3.1500 1.1250 ;
        RECT 1.0950 0.8025 1.2000 1.1250 ;
        RECT 0.7950 0.9750 1.0950 1.1250 ;
        RECT 0.6750 0.8250 0.7950 1.1250 ;
        RECT 0.3750 0.9750 0.6750 1.1250 ;
        RECT 0.2550 0.8550 0.3750 1.1250 ;
        RECT 0.0000 0.9750 0.2550 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 3.0150 0.1725 3.0750 0.2325 ;
        RECT 3.0150 0.8175 3.0750 0.8775 ;
        RECT 2.9100 0.4950 2.9700 0.5550 ;
        RECT 2.8050 0.3150 2.8650 0.3750 ;
        RECT 2.8050 0.6750 2.8650 0.7350 ;
        RECT 2.7000 0.4950 2.7600 0.5550 ;
        RECT 2.5950 0.1500 2.6550 0.2100 ;
        RECT 2.5950 0.8325 2.6550 0.8925 ;
        RECT 2.4900 0.4950 2.5500 0.5550 ;
        RECT 2.3850 0.3150 2.4450 0.3750 ;
        RECT 2.3850 0.6750 2.4450 0.7350 ;
        RECT 2.2800 0.4950 2.3400 0.5550 ;
        RECT 2.1750 0.1500 2.2350 0.2100 ;
        RECT 2.1750 0.8325 2.2350 0.8925 ;
        RECT 2.0700 0.4950 2.1300 0.5550 ;
        RECT 1.9650 0.3150 2.0250 0.3750 ;
        RECT 1.9650 0.6825 2.0250 0.7425 ;
        RECT 1.8600 0.4950 1.9200 0.5550 ;
        RECT 1.7550 0.1500 1.8150 0.2100 ;
        RECT 1.7550 0.8325 1.8150 0.8925 ;
        RECT 1.6500 0.4950 1.7100 0.5550 ;
        RECT 1.5450 0.3150 1.6050 0.3750 ;
        RECT 1.5450 0.6825 1.6050 0.7425 ;
        RECT 1.4400 0.4950 1.5000 0.5550 ;
        RECT 1.3350 0.1575 1.3950 0.2175 ;
        RECT 1.3350 0.8325 1.3950 0.8925 ;
        RECT 1.1250 0.1575 1.1850 0.2175 ;
        RECT 1.1250 0.8325 1.1850 0.8925 ;
        RECT 1.0200 0.4875 1.0800 0.5475 ;
        RECT 0.9150 0.3150 0.9750 0.3750 ;
        RECT 0.9150 0.6600 0.9750 0.7200 ;
        RECT 0.8100 0.4875 0.8700 0.5475 ;
        RECT 0.7050 0.1500 0.7650 0.2100 ;
        RECT 0.7050 0.8325 0.7650 0.8925 ;
        RECT 0.6000 0.4875 0.6600 0.5475 ;
        RECT 0.4950 0.3000 0.5550 0.3600 ;
        RECT 0.4950 0.6900 0.5550 0.7500 ;
        RECT 0.3900 0.4875 0.4500 0.5475 ;
        RECT 0.2850 0.1275 0.3450 0.1875 ;
        RECT 0.2850 0.8550 0.3450 0.9150 ;
        RECT 0.1800 0.4800 0.2400 0.5400 ;
        RECT 0.0750 0.2475 0.1350 0.3075 ;
        RECT 0.0750 0.7350 0.1350 0.7950 ;
        LAYER M1 ;
        RECT 2.9925 0.7950 3.0975 0.9000 ;
        RECT 1.3050 0.8250 2.9925 0.9000 ;
        RECT 2.3550 0.6525 2.8950 0.7500 ;
        RECT 0.5625 0.2925 2.8875 0.3975 ;
        RECT 1.4175 0.4725 2.1525 0.5775 ;
        RECT 1.3425 0.6750 2.0550 0.7500 ;
        RECT 1.2600 0.6525 1.3425 0.7500 ;
        RECT 0.5625 0.6525 1.2600 0.7275 ;
        RECT 0.4050 0.4800 1.1100 0.5550 ;
        RECT 0.4875 0.2625 0.5625 0.3975 ;
        RECT 0.4875 0.6525 0.5625 0.7875 ;
        RECT 0.3300 0.2625 0.4050 0.7800 ;
        RECT 0.1425 0.2625 0.3300 0.3375 ;
        RECT 0.1425 0.7050 0.3300 0.7800 ;
        RECT 0.0900 0.4125 0.2550 0.6225 ;
        RECT 0.0675 0.2175 0.1425 0.3375 ;
        RECT 0.0675 0.7050 0.1425 0.8250 ;
    END
END INR3_0111


MACRO INR3_1000
    CLASS CORE ;
    FOREIGN INR3_1000 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.0500 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.9975 0.3075 1.0125 0.9000 ;
        RECT 0.9375 0.1500 0.9975 0.9000 ;
        RECT 0.8925 0.1500 0.9375 0.3825 ;
        RECT 0.8850 0.7950 0.9375 0.9000 ;
        RECT 0.5625 0.3075 0.8925 0.3825 ;
        RECT 0.4875 0.1800 0.5625 0.3825 ;
        END
    END ZN
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.4575 0.5625 0.9225 0.6375 ;
        VIA 0.8100 0.6000 VIA12_square ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.2325 0.7125 0.6975 0.7875 ;
        VIA 0.5250 0.7500 VIA12_square ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.0975 0.4125 0.5625 0.4875 ;
        VIA 0.1800 0.4500 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.7950 -0.0750 1.0500 0.0750 ;
        RECT 0.6750 -0.0750 0.7950 0.2325 ;
        RECT 0.3750 -0.0750 0.6750 0.0750 ;
        RECT 0.2550 -0.0750 0.3750 0.1875 ;
        RECT 0.0000 -0.0750 0.2550 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.3750 0.9750 1.0500 1.1250 ;
        RECT 0.2550 0.8325 0.3750 1.1250 ;
        RECT 0.0000 0.9750 0.2550 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 0.9150 0.1725 0.9750 0.2325 ;
        RECT 0.9150 0.8175 0.9750 0.8775 ;
        RECT 0.8025 0.4950 0.8625 0.5550 ;
        RECT 0.7050 0.1575 0.7650 0.2175 ;
        RECT 0.5925 0.4950 0.6525 0.5550 ;
        RECT 0.4950 0.2100 0.5550 0.2700 ;
        RECT 0.3825 0.4875 0.4425 0.5475 ;
        RECT 0.2850 0.1200 0.3450 0.1800 ;
        RECT 0.2850 0.8400 0.3450 0.9000 ;
        RECT 0.1800 0.4875 0.2400 0.5475 ;
        RECT 0.0750 0.1725 0.1350 0.2325 ;
        RECT 0.0750 0.8175 0.1350 0.8775 ;
        LAYER M1 ;
        RECT 0.8025 0.4575 0.8625 0.7125 ;
        RECT 0.7575 0.4575 0.8025 0.8325 ;
        RECT 0.7275 0.6375 0.7575 0.8325 ;
        RECT 0.5625 0.4575 0.6525 0.7125 ;
        RECT 0.5475 0.4575 0.5625 0.8325 ;
        RECT 0.4875 0.6375 0.5475 0.8325 ;
        RECT 0.4125 0.4575 0.4425 0.5775 ;
        RECT 0.3375 0.2625 0.4125 0.7575 ;
        RECT 0.1575 0.2625 0.3375 0.3375 ;
        RECT 0.1575 0.6825 0.3375 0.7575 ;
        RECT 0.0975 0.4125 0.2625 0.6075 ;
        RECT 0.0525 0.1500 0.1575 0.3375 ;
        RECT 0.0525 0.6825 0.1575 0.9000 ;
    END
END INR3_1000


MACRO INR3_1010
    CLASS CORE ;
    FOREIGN INR3_1010 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.6800 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 1.1475 0.2625 1.6125 0.3375 ;
        RECT 1.0725 0.1650 1.1475 0.7950 ;
        RECT 0.9975 0.1650 1.0725 0.2550 ;
        RECT 0.8475 0.1500 0.9975 0.2550 ;
        VIA 1.4175 0.3000 VIA12_square ;
        VIA 1.1100 0.7125 VIA12_square ;
        VIA 0.9225 0.2025 VIA12_square ;
        END
    END ZN
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.7800 0.7125 0.9375 0.7875 ;
        RECT 0.6750 0.6225 0.7800 0.7875 ;
        RECT 0.3675 0.7125 0.6750 0.7875 ;
        VIA 0.7275 0.7050 VIA12_square ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.4350 0.4125 0.9000 0.4875 ;
        VIA 0.6150 0.4500 VIA12_square ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.0675 0.5625 0.5325 0.6375 ;
        VIA 0.2100 0.6000 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.6200 -0.0750 1.6800 0.0750 ;
        RECT 1.5450 -0.0750 1.6200 0.3075 ;
        RECT 1.1925 -0.0750 1.5450 0.0750 ;
        RECT 1.1100 -0.0750 1.1925 0.2100 ;
        RECT 0.1650 -0.0750 1.1100 0.0750 ;
        RECT 0.0450 -0.0750 0.1650 0.3150 ;
        RECT 0.0000 -0.0750 0.0450 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.6275 0.9750 1.6800 1.1250 ;
        RECT 1.5225 0.6450 1.6275 1.1250 ;
        RECT 0.3750 0.9750 1.5225 1.1250 ;
        RECT 0.2550 0.8700 0.3750 1.1250 ;
        RECT 0.0000 0.9750 0.2550 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.5450 0.2025 1.6050 0.2625 ;
        RECT 1.5450 0.6675 1.6050 0.7275 ;
        RECT 1.5450 0.8325 1.6050 0.8925 ;
        RECT 1.4400 0.4875 1.5000 0.5475 ;
        RECT 1.3350 0.1650 1.3950 0.2250 ;
        RECT 1.2300 0.4800 1.2900 0.5400 ;
        RECT 1.1250 0.1200 1.1850 0.1800 ;
        RECT 1.0200 0.4950 1.0800 0.5550 ;
        RECT 0.9150 0.1725 0.9750 0.2325 ;
        RECT 0.9150 0.6750 0.9750 0.7350 ;
        RECT 0.8100 0.4950 0.8700 0.5550 ;
        RECT 0.6000 0.4725 0.6600 0.5325 ;
        RECT 0.3900 0.4950 0.4500 0.5550 ;
        RECT 0.2850 0.2400 0.3450 0.3000 ;
        RECT 0.2850 0.8700 0.3450 0.9300 ;
        RECT 0.1800 0.4950 0.2400 0.5550 ;
        RECT 0.0750 0.2250 0.1350 0.2850 ;
        RECT 0.0750 0.7500 0.1350 0.8100 ;
        LAYER M1 ;
        RECT 1.4400 0.4725 1.5300 0.5625 ;
        RECT 1.3650 0.1500 1.4700 0.3975 ;
        RECT 1.3650 0.4725 1.4400 0.9000 ;
        RECT 1.2975 0.1500 1.3650 0.2400 ;
        RECT 0.5400 0.8250 1.3650 0.9000 ;
        RECT 1.1850 0.3150 1.2900 0.5700 ;
        RECT 1.0125 0.6750 1.2600 0.7500 ;
        RECT 0.6600 0.3150 1.1850 0.3900 ;
        RECT 0.8100 0.4650 1.1100 0.5700 ;
        RECT 0.8850 0.6450 1.0125 0.7500 ;
        RECT 0.6375 0.1500 1.0050 0.2400 ;
        RECT 0.7350 0.4650 0.8100 0.7425 ;
        RECT 0.6450 0.6675 0.7350 0.7425 ;
        RECT 0.5775 0.3150 0.6600 0.5625 ;
        RECT 0.4650 0.7200 0.5400 0.9000 ;
        RECT 0.4575 0.7200 0.4650 0.7950 ;
        RECT 0.3825 0.3000 0.4575 0.7950 ;
        RECT 0.3525 0.3000 0.3825 0.3750 ;
        RECT 0.1425 0.7200 0.3825 0.7950 ;
        RECT 0.2775 0.2100 0.3525 0.3750 ;
        RECT 0.1275 0.4500 0.2925 0.6450 ;
        RECT 0.0675 0.7200 0.1425 0.8400 ;
    END
END INR3_1010


MACRO INR4_0011
    CLASS CORE ;
    FOREIGN INR4_0011 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.9400 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 2.8275 0.3150 2.9025 0.8325 ;
        RECT 2.6625 0.3150 2.8275 0.3900 ;
        RECT 2.7975 0.6675 2.8275 0.8325 ;
        RECT 2.3400 0.6675 2.7975 0.7425 ;
        RECT 2.5875 0.2175 2.6625 0.3900 ;
        RECT 1.8225 0.3150 2.5875 0.3900 ;
        RECT 1.7475 0.2175 1.8225 0.3900 ;
        RECT 1.4025 0.3150 1.7475 0.3900 ;
        RECT 1.3275 0.2175 1.4025 0.3900 ;
        RECT 0.5625 0.3150 1.3275 0.3900 ;
        RECT 0.4875 0.2175 0.5625 0.3900 ;
        END
    END ZN
    PIN B3
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 2.4075 0.4500 2.5125 0.6375 ;
        RECT 1.9425 0.5625 2.4075 0.6375 ;
        VIA 2.4600 0.5250 VIA12_square ;
        END
    END B3
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.7475 0.4425 1.8225 0.7875 ;
        RECT 1.2825 0.7125 1.7475 0.7875 ;
        VIA 1.7850 0.5250 VIA12_square ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.3275 0.4425 1.4025 0.6375 ;
        RECT 0.8625 0.5625 1.3275 0.6375 ;
        VIA 1.3650 0.5250 VIA12_square ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.0900 0.4125 0.2550 0.6375 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 2.8950 -0.0750 2.9400 0.0750 ;
        RECT 2.7750 -0.0750 2.8950 0.2325 ;
        RECT 2.4750 -0.0750 2.7750 0.0750 ;
        RECT 2.3550 -0.0750 2.4750 0.2250 ;
        RECT 2.0550 -0.0750 2.3550 0.0750 ;
        RECT 1.9350 -0.0750 2.0550 0.2250 ;
        RECT 1.6350 -0.0750 1.9350 0.0750 ;
        RECT 1.5150 -0.0750 1.6350 0.2250 ;
        RECT 1.2150 -0.0750 1.5150 0.0750 ;
        RECT 1.0950 -0.0750 1.2150 0.2250 ;
        RECT 0.7950 -0.0750 1.0950 0.0750 ;
        RECT 0.6750 -0.0750 0.7950 0.2250 ;
        RECT 0.3750 -0.0750 0.6750 0.0750 ;
        RECT 0.2550 -0.0750 0.3750 0.1875 ;
        RECT 0.0000 -0.0750 0.2550 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.7950 0.9750 2.9400 1.1250 ;
        RECT 0.6750 0.8250 0.7950 1.1250 ;
        RECT 0.3750 0.9750 0.6750 1.1250 ;
        RECT 0.2550 0.8625 0.3750 1.1250 ;
        RECT 0.0000 0.9750 0.2550 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 2.8050 0.1725 2.8650 0.2325 ;
        RECT 2.8050 0.6825 2.8650 0.7425 ;
        RECT 2.6925 0.4950 2.7525 0.5550 ;
        RECT 2.5950 0.2475 2.6550 0.3075 ;
        RECT 2.5950 0.8325 2.6550 0.8925 ;
        RECT 2.4900 0.4950 2.5500 0.5550 ;
        RECT 2.3850 0.1575 2.4450 0.2175 ;
        RECT 2.3850 0.6750 2.4450 0.7350 ;
        RECT 2.2800 0.4950 2.3400 0.5550 ;
        RECT 2.1750 0.8250 2.2350 0.8850 ;
        RECT 2.0700 0.4950 2.1300 0.5550 ;
        RECT 1.9650 0.1575 2.0250 0.2175 ;
        RECT 1.9650 0.6825 2.0250 0.7425 ;
        RECT 1.8600 0.4950 1.9200 0.5550 ;
        RECT 1.7550 0.2475 1.8150 0.3075 ;
        RECT 1.7550 0.8250 1.8150 0.8850 ;
        RECT 1.6500 0.4950 1.7100 0.5550 ;
        RECT 1.5450 0.1575 1.6050 0.2175 ;
        RECT 1.5450 0.7500 1.6050 0.8100 ;
        RECT 1.4400 0.4950 1.5000 0.5550 ;
        RECT 1.3350 0.2475 1.3950 0.3075 ;
        RECT 1.3350 0.6825 1.3950 0.7425 ;
        RECT 1.2300 0.4950 1.2900 0.5550 ;
        RECT 1.1250 0.1575 1.1850 0.2175 ;
        RECT 1.1250 0.8325 1.1850 0.8925 ;
        RECT 1.0275 0.4950 1.0875 0.5550 ;
        RECT 0.9150 0.6825 0.9750 0.7425 ;
        RECT 0.8025 0.4950 0.8625 0.5550 ;
        RECT 0.7050 0.1575 0.7650 0.2175 ;
        RECT 0.7050 0.8325 0.7650 0.8925 ;
        RECT 0.6000 0.4950 0.6600 0.5550 ;
        RECT 0.4950 0.2475 0.5550 0.3075 ;
        RECT 0.4950 0.7200 0.5550 0.7800 ;
        RECT 0.3900 0.4950 0.4500 0.5550 ;
        RECT 0.2850 0.1275 0.3450 0.1875 ;
        RECT 0.2850 0.8625 0.3450 0.9225 ;
        RECT 0.1800 0.4800 0.2400 0.5400 ;
        RECT 0.0750 0.2475 0.1350 0.3075 ;
        RECT 0.0750 0.7425 0.1350 0.8025 ;
        LAYER M1 ;
        RECT 2.2800 0.4650 2.7525 0.5850 ;
        RECT 1.8450 0.8250 2.6850 0.9000 ;
        RECT 1.7325 0.4725 2.1600 0.5625 ;
        RECT 1.9350 0.6450 2.0550 0.7500 ;
        RECT 1.6125 0.6600 1.9350 0.7350 ;
        RECT 1.7250 0.8100 1.8450 0.9000 ;
        RECT 1.6125 0.4725 1.7325 0.5775 ;
        RECT 1.5375 0.6600 1.6125 0.9000 ;
        RECT 1.0950 0.8250 1.5375 0.9000 ;
        RECT 0.9975 0.4725 1.5225 0.5775 ;
        RECT 0.5625 0.6750 1.4250 0.7500 ;
        RECT 0.4050 0.4875 0.8925 0.5625 ;
        RECT 0.4875 0.6750 0.5625 0.8100 ;
        RECT 0.3300 0.2625 0.4050 0.7875 ;
        RECT 0.1425 0.2625 0.3300 0.3375 ;
        RECT 0.1425 0.7125 0.3300 0.7875 ;
        RECT 0.0675 0.2175 0.1425 0.3375 ;
        RECT 0.0675 0.7125 0.1425 0.8325 ;
    END
END INR4_0011


MACRO INR4_0111
    CLASS CORE ;
    FOREIGN INR4_0111 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.2000 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 3.5175 0.2625 3.8325 0.7875 ;
        VIA 3.6750 0.3450 VIA12_slot ;
        VIA 3.6750 0.7050 VIA12_slot ;
        END
    END ZN
    PIN B3
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 3.2550 0.4425 3.3300 0.6375 ;
        RECT 2.7900 0.5625 3.2550 0.6375 ;
        VIA 3.2925 0.5250 VIA12_square ;
        END
    END B3
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 2.3775 0.4500 2.4525 0.6375 ;
        RECT 1.9125 0.5625 2.3775 0.6375 ;
        VIA 2.4150 0.5400 VIA12_square ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.5375 0.4500 1.6125 0.6375 ;
        RECT 1.0725 0.5625 1.5375 0.6375 ;
        VIA 1.5750 0.5400 VIA12_square ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.0900 0.4125 0.5550 0.4875 ;
        VIA 0.1725 0.4500 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 4.1325 -0.0750 4.2000 0.0750 ;
        RECT 4.0575 -0.0750 4.1325 0.2625 ;
        RECT 3.7350 -0.0750 4.0575 0.0750 ;
        RECT 3.6150 -0.0750 3.7350 0.2175 ;
        RECT 3.3150 -0.0750 3.6150 0.0750 ;
        RECT 3.1950 -0.0750 3.3150 0.2175 ;
        RECT 3.1050 -0.0750 3.1950 0.0750 ;
        RECT 2.9850 -0.0750 3.1050 0.2175 ;
        RECT 2.6850 -0.0750 2.9850 0.0750 ;
        RECT 2.5650 -0.0750 2.6850 0.2175 ;
        RECT 2.2650 -0.0750 2.5650 0.0750 ;
        RECT 2.1450 -0.0750 2.2650 0.2175 ;
        RECT 1.8450 -0.0750 2.1450 0.0750 ;
        RECT 1.7250 -0.0750 1.8450 0.2175 ;
        RECT 1.4250 -0.0750 1.7250 0.0750 ;
        RECT 1.3050 -0.0750 1.4250 0.2175 ;
        RECT 1.2150 -0.0750 1.3050 0.0750 ;
        RECT 1.0950 -0.0750 1.2150 0.2175 ;
        RECT 0.7950 -0.0750 1.0950 0.0750 ;
        RECT 0.6750 -0.0750 0.7950 0.2175 ;
        RECT 0.3750 -0.0750 0.6750 0.0750 ;
        RECT 0.2550 -0.0750 0.3750 0.1875 ;
        RECT 0.0000 -0.0750 0.2550 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.2000 0.9750 4.2000 1.1250 ;
        RECT 1.0950 0.8025 1.2000 1.1250 ;
        RECT 0.7875 0.9750 1.0950 1.1250 ;
        RECT 0.6825 0.8100 0.7875 1.1250 ;
        RECT 0.3750 0.9750 0.6825 1.1250 ;
        RECT 0.2550 0.8550 0.3750 1.1250 ;
        RECT 0.0000 0.9750 0.2550 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 4.0650 0.1725 4.1250 0.2325 ;
        RECT 4.0650 0.8175 4.1250 0.8775 ;
        RECT 3.9600 0.4950 4.0200 0.5550 ;
        RECT 3.8550 0.3150 3.9150 0.3750 ;
        RECT 3.8550 0.6675 3.9150 0.7275 ;
        RECT 3.7500 0.4950 3.8100 0.5550 ;
        RECT 3.6450 0.1500 3.7050 0.2100 ;
        RECT 3.6450 0.8325 3.7050 0.8925 ;
        RECT 3.5400 0.4950 3.6000 0.5550 ;
        RECT 3.4350 0.3150 3.4950 0.3750 ;
        RECT 3.4350 0.6675 3.4950 0.7275 ;
        RECT 3.3300 0.4950 3.3900 0.5550 ;
        RECT 3.2250 0.1575 3.2850 0.2175 ;
        RECT 3.2250 0.7575 3.2850 0.8175 ;
        RECT 3.0150 0.1575 3.0750 0.2175 ;
        RECT 3.0150 0.8325 3.0750 0.8925 ;
        RECT 2.9100 0.4950 2.9700 0.5550 ;
        RECT 2.8050 0.3150 2.8650 0.3750 ;
        RECT 2.8050 0.6825 2.8650 0.7425 ;
        RECT 2.7000 0.4950 2.7600 0.5550 ;
        RECT 2.5950 0.1500 2.6550 0.2100 ;
        RECT 2.5950 0.8325 2.6550 0.8925 ;
        RECT 2.4900 0.4950 2.5500 0.5550 ;
        RECT 2.3850 0.3150 2.4450 0.3750 ;
        RECT 2.3850 0.6825 2.4450 0.7425 ;
        RECT 2.2800 0.4950 2.3400 0.5550 ;
        RECT 2.1750 0.1500 2.2350 0.2100 ;
        RECT 2.1750 0.8325 2.2350 0.8925 ;
        RECT 2.0700 0.4950 2.1300 0.5550 ;
        RECT 1.9650 0.3150 2.0250 0.3750 ;
        RECT 1.9650 0.6825 2.0250 0.7425 ;
        RECT 1.8600 0.4950 1.9200 0.5550 ;
        RECT 1.7550 0.1500 1.8150 0.2100 ;
        RECT 1.7550 0.8325 1.8150 0.8925 ;
        RECT 1.6500 0.4950 1.7100 0.5550 ;
        RECT 1.5450 0.3150 1.6050 0.3750 ;
        RECT 1.5450 0.6825 1.6050 0.7425 ;
        RECT 1.4400 0.4950 1.5000 0.5550 ;
        RECT 1.3350 0.1575 1.3950 0.2175 ;
        RECT 1.3350 0.8325 1.3950 0.8925 ;
        RECT 1.1250 0.1575 1.1850 0.2175 ;
        RECT 1.1250 0.8325 1.1850 0.8925 ;
        RECT 1.0200 0.4950 1.0800 0.5550 ;
        RECT 0.9150 0.3150 0.9750 0.3750 ;
        RECT 0.9150 0.6675 0.9750 0.7275 ;
        RECT 0.8100 0.4950 0.8700 0.5550 ;
        RECT 0.7050 0.1500 0.7650 0.2100 ;
        RECT 0.7050 0.8325 0.7650 0.8925 ;
        RECT 0.6000 0.4950 0.6600 0.5550 ;
        RECT 0.4950 0.2925 0.5550 0.3525 ;
        RECT 0.4950 0.6825 0.5550 0.7425 ;
        RECT 0.3900 0.4950 0.4500 0.5550 ;
        RECT 0.2850 0.1275 0.3450 0.1875 ;
        RECT 0.2850 0.8550 0.3450 0.9150 ;
        RECT 0.1800 0.4800 0.2400 0.5400 ;
        RECT 0.0750 0.2475 0.1350 0.3075 ;
        RECT 0.0750 0.7350 0.1350 0.7950 ;
        LAYER M1 ;
        RECT 4.0425 0.7875 4.1475 0.9000 ;
        RECT 3.2100 0.4875 4.0650 0.5625 ;
        RECT 3.2925 0.8250 4.0425 0.9000 ;
        RECT 0.5625 0.2925 3.9450 0.3975 ;
        RECT 3.4125 0.6450 3.9375 0.7500 ;
        RECT 3.2175 0.6750 3.2925 0.9000 ;
        RECT 2.3550 0.6750 3.2175 0.7500 ;
        RECT 1.3050 0.8250 3.1050 0.9000 ;
        RECT 2.2575 0.4725 2.9925 0.5775 ;
        RECT 1.4175 0.4725 2.1525 0.5775 ;
        RECT 1.3425 0.6750 2.0550 0.7500 ;
        RECT 1.2600 0.6525 1.3425 0.7500 ;
        RECT 0.5625 0.6525 1.2600 0.7275 ;
        RECT 0.4050 0.4875 1.1100 0.5625 ;
        RECT 0.4875 0.2400 0.5625 0.3975 ;
        RECT 0.4875 0.6525 0.5625 0.7875 ;
        RECT 0.3300 0.2625 0.4050 0.7800 ;
        RECT 0.1425 0.2625 0.3300 0.3375 ;
        RECT 0.1425 0.7050 0.3300 0.7800 ;
        RECT 0.0900 0.4125 0.2550 0.6300 ;
        RECT 0.0675 0.2175 0.1425 0.3375 ;
        RECT 0.0675 0.7050 0.1425 0.8250 ;
    END
END INR4_0111


MACRO INR4_1000
    CLASS CORE ;
    FOREIGN INR4_1000 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.2600 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 1.1475 0.3075 1.2225 0.9000 ;
        RECT 0.9825 0.3075 1.1475 0.3825 ;
        RECT 1.1025 0.7950 1.1475 0.9000 ;
        RECT 0.9075 0.1800 0.9825 0.3825 ;
        RECT 0.5625 0.3075 0.9075 0.3825 ;
        RECT 0.4875 0.1800 0.5625 0.3825 ;
        END
    END ZN
    PIN B3
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.7275 0.7125 1.1925 0.7875 ;
        VIA 0.9825 0.7500 VIA12_square ;
        END
    END B3
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.4350 0.5625 0.9000 0.6375 ;
        VIA 0.7800 0.6000 VIA12_square ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.1425 0.7125 0.6075 0.7875 ;
        VIA 0.5250 0.7500 VIA12_square ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.0900 0.4125 0.5550 0.4875 ;
        VIA 0.1725 0.4500 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.2150 -0.0750 1.2600 0.0750 ;
        RECT 1.0950 -0.0750 1.2150 0.2175 ;
        RECT 0.7950 -0.0750 1.0950 0.0750 ;
        RECT 0.6750 -0.0750 0.7950 0.2100 ;
        RECT 0.3750 -0.0750 0.6750 0.0750 ;
        RECT 0.2550 -0.0750 0.3750 0.1875 ;
        RECT 0.0000 -0.0750 0.2550 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.3750 0.9750 1.2600 1.1250 ;
        RECT 0.2550 0.8475 0.3750 1.1250 ;
        RECT 0.0000 0.9750 0.2550 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.1250 0.1575 1.1850 0.2175 ;
        RECT 1.1250 0.8175 1.1850 0.8775 ;
        RECT 1.0125 0.5100 1.0725 0.5700 ;
        RECT 0.9150 0.2100 0.9750 0.2700 ;
        RECT 0.8100 0.5175 0.8700 0.5775 ;
        RECT 0.7050 0.1200 0.7650 0.1800 ;
        RECT 0.6000 0.5250 0.6600 0.5850 ;
        RECT 0.4950 0.2100 0.5550 0.2700 ;
        RECT 0.3900 0.5100 0.4500 0.5700 ;
        RECT 0.2850 0.1200 0.3450 0.1800 ;
        RECT 0.2850 0.8625 0.3450 0.9225 ;
        RECT 0.1800 0.5100 0.2400 0.5700 ;
        RECT 0.0750 0.1725 0.1350 0.2325 ;
        RECT 0.0750 0.8175 0.1350 0.8775 ;
        LAYER M1 ;
        RECT 1.0200 0.4575 1.0725 0.6000 ;
        RECT 0.9450 0.4575 1.0200 0.8325 ;
        RECT 0.8325 0.4575 0.8700 0.6075 ;
        RECT 0.7425 0.4575 0.8325 0.7725 ;
        RECT 0.5775 0.4875 0.6675 0.8325 ;
        RECT 0.4875 0.6675 0.5775 0.8325 ;
        RECT 0.4125 0.4875 0.4725 0.5925 ;
        RECT 0.3375 0.2625 0.4125 0.7725 ;
        RECT 0.1575 0.2625 0.3375 0.3375 ;
        RECT 0.1575 0.6975 0.3375 0.7725 ;
        RECT 0.0900 0.4125 0.2550 0.6225 ;
        RECT 0.0525 0.1500 0.1575 0.3375 ;
        RECT 0.0525 0.6975 0.1575 0.9000 ;
    END
END INR4_1000


MACRO INR4_1010
    CLASS CORE ;
    FOREIGN INR4_1010 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.3100 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 1.8225 0.1425 1.9275 0.3375 ;
        RECT 1.3125 0.2625 1.8225 0.3375 ;
        RECT 1.3125 0.6600 1.4325 0.7350 ;
        RECT 1.2375 0.1950 1.3125 0.7350 ;
        RECT 0.6525 0.1950 1.2375 0.2700 ;
        VIA 1.8750 0.2250 VIA12_square ;
        VIA 1.3500 0.6975 VIA12_square ;
        VIA 0.7350 0.2325 VIA12_square ;
        END
    END ZN
    PIN B3
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.4925 0.4125 1.9575 0.4875 ;
        VIA 1.7325 0.4500 VIA12_square ;
        END
    END B3
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 2.1675 0.3675 2.2425 0.5400 ;
        RECT 2.0850 0.4650 2.1675 0.5400 ;
        RECT 2.0100 0.4650 2.0850 0.7350 ;
        RECT 1.5750 0.6600 2.0100 0.7350 ;
        RECT 1.5000 0.4200 1.5750 0.7350 ;
        RECT 1.4325 0.4200 1.5000 0.5400 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.3900 0.5625 0.8550 0.6375 ;
        VIA 0.6600 0.6000 VIA12_square ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1425 0.4350 0.2400 0.5550 ;
        RECT 0.0675 0.3675 0.1425 0.6825 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 2.2650 -0.0750 2.3100 0.0750 ;
        RECT 2.1450 -0.0750 2.2650 0.2625 ;
        RECT 1.6350 -0.0750 2.1450 0.0750 ;
        RECT 1.5150 -0.0750 1.6350 0.2475 ;
        RECT 0.9900 -0.0750 1.5150 0.0750 ;
        RECT 0.9000 -0.0750 0.9900 0.3075 ;
        RECT 0.5850 -0.0750 0.9000 0.0750 ;
        RECT 0.4650 -0.0750 0.5850 0.2400 ;
        RECT 0.1650 -0.0750 0.4650 0.0750 ;
        RECT 0.0450 -0.0750 0.1650 0.2625 ;
        RECT 0.0000 -0.0750 0.0450 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.0125 0.9750 2.3100 1.1250 ;
        RECT 0.9075 0.8100 1.0125 1.1250 ;
        RECT 0.1650 0.9750 0.9075 1.1250 ;
        RECT 0.0450 0.7875 0.1650 1.1250 ;
        RECT 0.0000 0.9750 0.0450 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 2.1750 0.1725 2.2350 0.2325 ;
        RECT 2.1750 0.8325 2.2350 0.8925 ;
        RECT 2.0700 0.4725 2.1300 0.5325 ;
        RECT 1.9650 0.1875 2.0250 0.2475 ;
        RECT 1.8600 0.4950 1.9200 0.5550 ;
        RECT 1.7550 0.1875 1.8150 0.2475 ;
        RECT 1.7550 0.8175 1.8150 0.8775 ;
        RECT 1.6500 0.4950 1.7100 0.5550 ;
        RECT 1.5450 0.1575 1.6050 0.2175 ;
        RECT 1.4400 0.4500 1.5000 0.5100 ;
        RECT 1.2300 0.3750 1.2900 0.4350 ;
        RECT 1.0200 0.4950 1.0800 0.5550 ;
        RECT 0.9150 0.2100 0.9750 0.2700 ;
        RECT 0.9150 0.8400 0.9750 0.9000 ;
        RECT 0.8100 0.4950 0.8700 0.5550 ;
        RECT 0.7050 0.2025 0.7650 0.2625 ;
        RECT 0.6000 0.4950 0.6600 0.5550 ;
        RECT 0.4950 0.1575 0.5550 0.2175 ;
        RECT 0.4950 0.8250 0.5550 0.8850 ;
        RECT 0.2850 0.2400 0.3450 0.3000 ;
        RECT 0.2850 0.6750 0.3450 0.7350 ;
        RECT 0.1800 0.4650 0.2400 0.5250 ;
        RECT 0.0750 0.1725 0.1350 0.2325 ;
        RECT 0.0750 0.8325 0.1350 0.8925 ;
        LAYER M1 ;
        RECT 2.1600 0.7800 2.2650 0.9000 ;
        RECT 1.9500 0.8100 2.1600 0.9000 ;
        RECT 1.7250 0.1725 2.0550 0.2775 ;
        RECT 1.8150 0.4650 1.9200 0.5850 ;
        RECT 1.4175 0.8100 1.8450 0.8850 ;
        RECT 1.6500 0.4125 1.8150 0.5850 ;
        RECT 1.3125 0.6150 1.4175 0.8850 ;
        RECT 1.2300 0.3450 1.2975 0.4650 ;
        RECT 1.1550 0.3450 1.2300 0.7350 ;
        RECT 0.6975 0.6600 1.1550 0.7350 ;
        RECT 0.8100 0.4650 1.0800 0.5850 ;
        RECT 0.6600 0.1500 0.8100 0.3600 ;
        RECT 0.4500 0.8100 0.8025 0.9000 ;
        RECT 0.6225 0.4950 0.6975 0.7350 ;
        RECT 0.5475 0.4950 0.6225 0.6075 ;
        RECT 0.3900 0.3150 0.5550 0.4200 ;
        RECT 0.3150 0.2100 0.3900 0.7650 ;
        RECT 0.2775 0.2100 0.3150 0.3300 ;
        RECT 0.2775 0.6450 0.3150 0.7650 ;
        LAYER VIA1 ;
        RECT 1.9950 0.8100 2.0700 0.8850 ;
        RECT 0.9600 0.4800 1.0350 0.5550 ;
        RECT 0.6600 0.8100 0.7350 0.8850 ;
        RECT 0.4350 0.3450 0.5100 0.4200 ;
        LAYER M2 ;
        RECT 0.6150 0.8100 2.2050 0.8850 ;
        RECT 0.9600 0.3450 1.0350 0.6000 ;
        RECT 0.3900 0.3450 0.9600 0.4200 ;
    END
END INR4_1010


MACRO INV_0001
    CLASS CORE ;
    FOREIGN INV_0001 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.8400 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.7275 0.2025 0.8025 0.8400 ;
        RECT 0.6975 0.2025 0.7275 0.3750 ;
        RECT 0.6975 0.6525 0.7275 0.8400 ;
        RECT 0.3525 0.3000 0.6975 0.3750 ;
        RECT 0.3525 0.6525 0.6975 0.7275 ;
        RECT 0.2775 0.2025 0.3525 0.3750 ;
        RECT 0.2775 0.6525 0.3525 0.8400 ;
        END
    END ZN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1425 0.4500 0.6525 0.5700 ;
        RECT 0.0675 0.3675 0.1425 0.6825 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.5850 -0.0750 0.8400 0.0750 ;
        RECT 0.4650 -0.0750 0.5850 0.2250 ;
        RECT 0.1425 -0.0750 0.4650 0.0750 ;
        RECT 0.0675 -0.0750 0.1425 0.2475 ;
        RECT 0.0000 -0.0750 0.0675 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.5850 0.9750 0.8400 1.1250 ;
        RECT 0.4650 0.8175 0.5850 1.1250 ;
        RECT 0.1425 0.9750 0.4650 1.1250 ;
        RECT 0.0675 0.8025 0.1425 1.1250 ;
        RECT 0.0000 0.9750 0.0675 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 0.7050 0.2325 0.7650 0.2925 ;
        RECT 0.7050 0.7500 0.7650 0.8100 ;
        RECT 0.5925 0.4800 0.6525 0.5400 ;
        RECT 0.4950 0.1500 0.5550 0.2100 ;
        RECT 0.4950 0.8325 0.5550 0.8925 ;
        RECT 0.3900 0.4800 0.4500 0.5400 ;
        RECT 0.2850 0.2325 0.3450 0.2925 ;
        RECT 0.2850 0.7500 0.3450 0.8100 ;
        RECT 0.1800 0.4800 0.2400 0.5400 ;
        RECT 0.0750 0.1575 0.1350 0.2175 ;
        RECT 0.0750 0.8325 0.1350 0.8925 ;
    END
END INV_0001


MACRO INV_0011
    CLASS CORE ;
    FOREIGN INV_0011 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.6300 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.5175 0.3075 0.5925 0.7275 ;
        RECT 0.3525 0.3075 0.5175 0.3825 ;
        RECT 0.3525 0.6525 0.5175 0.7275 ;
        RECT 0.2775 0.2175 0.3525 0.3825 ;
        RECT 0.2775 0.6525 0.3525 0.8325 ;
        END
    END ZN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1425 0.4575 0.4425 0.5775 ;
        RECT 0.0675 0.3675 0.1425 0.6825 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.5850 -0.0750 0.6300 0.0750 ;
        RECT 0.4650 -0.0750 0.5850 0.2325 ;
        RECT 0.1425 -0.0750 0.4650 0.0750 ;
        RECT 0.0675 -0.0750 0.1425 0.2475 ;
        RECT 0.0000 -0.0750 0.0675 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.5775 0.9750 0.6300 1.1250 ;
        RECT 0.4725 0.8025 0.5775 1.1250 ;
        RECT 0.1425 0.9750 0.4725 1.1250 ;
        RECT 0.0675 0.8025 0.1425 1.1250 ;
        RECT 0.0000 0.9750 0.0675 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 0.4950 0.1575 0.5550 0.2175 ;
        RECT 0.4950 0.8250 0.5550 0.8850 ;
        RECT 0.3825 0.4875 0.4425 0.5475 ;
        RECT 0.2850 0.2550 0.3450 0.3150 ;
        RECT 0.2850 0.7425 0.3450 0.8025 ;
        RECT 0.1800 0.4875 0.2400 0.5475 ;
        RECT 0.0750 0.1575 0.1350 0.2175 ;
        RECT 0.0750 0.8325 0.1350 0.8925 ;
    END
END INV_0011


MACRO INV_0100
    CLASS CORE ;
    FOREIGN INV_0100 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.8900 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 1.1025 0.2775 1.2600 0.3975 ;
        RECT 1.1025 0.6525 1.2600 0.7725 ;
        RECT 0.7875 0.2775 1.1025 0.7725 ;
        RECT 0.6300 0.2775 0.7875 0.3975 ;
        RECT 0.6300 0.6525 0.7875 0.7725 ;
        VIA 1.1025 0.3375 VIA12_slot ;
        VIA 1.1025 0.7125 VIA12_slot ;
        VIA 0.7875 0.3375 VIA12_slot ;
        VIA 0.7875 0.7125 VIA12_slot ;
        END
    END ZN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1425 0.4725 1.7850 0.5475 ;
        RECT 0.0675 0.3675 0.1425 0.6825 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.8450 -0.0750 1.8900 0.0750 ;
        RECT 1.7250 -0.0750 1.8450 0.2925 ;
        RECT 1.4250 -0.0750 1.7250 0.0750 ;
        RECT 1.3050 -0.0750 1.4250 0.2025 ;
        RECT 1.0050 -0.0750 1.3050 0.0750 ;
        RECT 0.8850 -0.0750 1.0050 0.2025 ;
        RECT 0.5850 -0.0750 0.8850 0.0750 ;
        RECT 0.4650 -0.0750 0.5850 0.2025 ;
        RECT 0.1425 -0.0750 0.4650 0.0750 ;
        RECT 0.0675 -0.0750 0.1425 0.2475 ;
        RECT 0.0000 -0.0750 0.0675 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.8450 0.9750 1.8900 1.1250 ;
        RECT 1.7250 0.6600 1.8450 1.1250 ;
        RECT 1.4250 0.9750 1.7250 1.1250 ;
        RECT 1.3050 0.8475 1.4250 1.1250 ;
        RECT 1.0050 0.9750 1.3050 1.1250 ;
        RECT 0.8850 0.8475 1.0050 1.1250 ;
        RECT 0.5850 0.9750 0.8850 1.1250 ;
        RECT 0.4650 0.8475 0.5850 1.1250 ;
        RECT 0.1425 0.9750 0.4650 1.1250 ;
        RECT 0.0675 0.8025 0.1425 1.1250 ;
        RECT 0.0000 0.9750 0.0675 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.7550 0.2175 1.8150 0.2775 ;
        RECT 1.7550 0.6675 1.8150 0.7275 ;
        RECT 1.7550 0.8325 1.8150 0.8925 ;
        RECT 1.6500 0.4800 1.7100 0.5400 ;
        RECT 1.5450 0.3075 1.6050 0.3675 ;
        RECT 1.5450 0.6825 1.6050 0.7425 ;
        RECT 1.4400 0.4800 1.5000 0.5400 ;
        RECT 1.3350 0.1350 1.3950 0.1950 ;
        RECT 1.3350 0.8550 1.3950 0.9150 ;
        RECT 1.2300 0.4800 1.2900 0.5400 ;
        RECT 1.1250 0.3075 1.1850 0.3675 ;
        RECT 1.1250 0.6825 1.1850 0.7425 ;
        RECT 1.0200 0.4800 1.0800 0.5400 ;
        RECT 0.9150 0.1350 0.9750 0.1950 ;
        RECT 0.9150 0.8550 0.9750 0.9150 ;
        RECT 0.8100 0.4800 0.8700 0.5400 ;
        RECT 0.7050 0.3075 0.7650 0.3675 ;
        RECT 0.7050 0.6825 0.7650 0.7425 ;
        RECT 0.6000 0.4800 0.6600 0.5400 ;
        RECT 0.4950 0.1350 0.5550 0.1950 ;
        RECT 0.4950 0.8550 0.5550 0.9150 ;
        RECT 0.3900 0.4800 0.4500 0.5400 ;
        RECT 0.2850 0.3075 0.3450 0.3675 ;
        RECT 0.2850 0.6825 0.3450 0.7425 ;
        RECT 0.1800 0.4800 0.2400 0.5400 ;
        RECT 0.0750 0.1575 0.1350 0.2175 ;
        RECT 0.0750 0.8325 0.1350 0.8925 ;
        LAYER M1 ;
        RECT 0.2775 0.2775 1.6200 0.3975 ;
        RECT 0.2775 0.6525 1.6200 0.7725 ;
        LAYER M2 ;
        RECT 0.6300 0.6525 0.7575 0.7725 ;
        RECT 1.1325 0.2775 1.2600 0.3975 ;
        RECT 1.1325 0.6525 1.2600 0.7725 ;
        RECT 0.6300 0.2775 0.7575 0.3975 ;
    END
END INV_0100


MACRO INV_0101
    CLASS CORE ;
    FOREIGN INV_0101 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.7300 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 1.5225 0.2775 1.6800 0.3975 ;
        RECT 1.5225 0.6525 1.6800 0.7725 ;
        RECT 1.2075 0.2775 1.5225 0.7725 ;
        RECT 1.0500 0.2775 1.2075 0.3975 ;
        RECT 1.0500 0.6525 1.2075 0.7725 ;
        VIA 1.5225 0.3375 VIA12_slot ;
        VIA 1.5225 0.7125 VIA12_slot ;
        VIA 1.2075 0.3375 VIA12_slot ;
        VIA 1.2075 0.7125 VIA12_slot ;
        END
    END ZN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1425 0.4725 2.6250 0.5475 ;
        RECT 0.0675 0.3675 0.1425 0.6825 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 2.6850 -0.0750 2.7300 0.0750 ;
        RECT 2.5650 -0.0750 2.6850 0.2925 ;
        RECT 2.2650 -0.0750 2.5650 0.0750 ;
        RECT 2.1450 -0.0750 2.2650 0.2025 ;
        RECT 1.8450 -0.0750 2.1450 0.0750 ;
        RECT 1.7250 -0.0750 1.8450 0.2025 ;
        RECT 1.4250 -0.0750 1.7250 0.0750 ;
        RECT 1.3050 -0.0750 1.4250 0.2025 ;
        RECT 1.0050 -0.0750 1.3050 0.0750 ;
        RECT 0.8850 -0.0750 1.0050 0.2025 ;
        RECT 0.5850 -0.0750 0.8850 0.0750 ;
        RECT 0.4650 -0.0750 0.5850 0.2025 ;
        RECT 0.1425 -0.0750 0.4650 0.0750 ;
        RECT 0.0675 -0.0750 0.1425 0.2475 ;
        RECT 0.0000 -0.0750 0.0675 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 2.6850 0.9750 2.7300 1.1250 ;
        RECT 2.5650 0.6600 2.6850 1.1250 ;
        RECT 2.2650 0.9750 2.5650 1.1250 ;
        RECT 2.1450 0.8475 2.2650 1.1250 ;
        RECT 1.8450 0.9750 2.1450 1.1250 ;
        RECT 1.7250 0.8475 1.8450 1.1250 ;
        RECT 1.4250 0.9750 1.7250 1.1250 ;
        RECT 1.3050 0.8475 1.4250 1.1250 ;
        RECT 1.0050 0.9750 1.3050 1.1250 ;
        RECT 0.8850 0.8475 1.0050 1.1250 ;
        RECT 0.5850 0.9750 0.8850 1.1250 ;
        RECT 0.4650 0.8475 0.5850 1.1250 ;
        RECT 0.1425 0.9750 0.4650 1.1250 ;
        RECT 0.0675 0.8025 0.1425 1.1250 ;
        RECT 0.0000 0.9750 0.0675 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 2.5950 0.2250 2.6550 0.2850 ;
        RECT 2.5950 0.6675 2.6550 0.7275 ;
        RECT 2.5950 0.8325 2.6550 0.8925 ;
        RECT 2.3850 0.6825 2.4450 0.7425 ;
        RECT 2.2800 0.4800 2.3400 0.5400 ;
        RECT 2.1750 0.1350 2.2350 0.1950 ;
        RECT 2.1750 0.8550 2.2350 0.9150 ;
        RECT 2.0700 0.4800 2.1300 0.5400 ;
        RECT 1.9650 0.3075 2.0250 0.3675 ;
        RECT 1.9650 0.6825 2.0250 0.7425 ;
        RECT 1.8600 0.4800 1.9200 0.5400 ;
        RECT 1.7550 0.1350 1.8150 0.1950 ;
        RECT 1.7550 0.8550 1.8150 0.9150 ;
        RECT 1.6500 0.4800 1.7100 0.5400 ;
        RECT 1.5450 0.3075 1.6050 0.3675 ;
        RECT 1.5450 0.6825 1.6050 0.7425 ;
        RECT 1.4400 0.4800 1.5000 0.5400 ;
        RECT 1.3350 0.1350 1.3950 0.1950 ;
        RECT 1.3350 0.8550 1.3950 0.9150 ;
        RECT 1.2300 0.4800 1.2900 0.5400 ;
        RECT 1.1250 0.3075 1.1850 0.3675 ;
        RECT 1.1250 0.6825 1.1850 0.7425 ;
        RECT 1.0200 0.4800 1.0800 0.5400 ;
        RECT 0.9150 0.1350 0.9750 0.1950 ;
        RECT 0.9150 0.8550 0.9750 0.9150 ;
        RECT 0.8100 0.4800 0.8700 0.5400 ;
        RECT 0.7050 0.3075 0.7650 0.3675 ;
        RECT 0.7050 0.6825 0.7650 0.7425 ;
        RECT 0.6000 0.4800 0.6600 0.5400 ;
        RECT 0.4950 0.1350 0.5550 0.1950 ;
        RECT 0.4950 0.8550 0.5550 0.9150 ;
        RECT 0.3900 0.4800 0.4500 0.5400 ;
        RECT 0.2850 0.3075 0.3450 0.3675 ;
        RECT 0.2850 0.6825 0.3450 0.7425 ;
        RECT 0.1800 0.4800 0.2400 0.5400 ;
        RECT 0.0750 0.1575 0.1350 0.2175 ;
        RECT 0.0750 0.8325 0.1350 0.8925 ;
        RECT 2.4900 0.4800 2.5500 0.5400 ;
        RECT 2.3850 0.3075 2.4450 0.3675 ;
        LAYER M1 ;
        RECT 0.2775 0.2775 2.4600 0.3975 ;
        RECT 0.2775 0.6525 2.4600 0.7725 ;
        LAYER M2 ;
        RECT 1.5525 0.2775 1.6800 0.3975 ;
        RECT 1.5525 0.6525 1.6800 0.7725 ;
        RECT 1.0500 0.2775 1.1775 0.3975 ;
        RECT 1.0500 0.6525 1.1775 0.7725 ;
    END
END INV_0101


MACRO INV_0110
    CLASS CORE ;
    FOREIGN INV_0110 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.4700 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 0.8925 0.2775 1.0500 0.3975 ;
        RECT 0.8925 0.6525 1.0500 0.7725 ;
        RECT 0.5775 0.2775 0.8925 0.7725 ;
        RECT 0.4200 0.2775 0.5775 0.3975 ;
        RECT 0.4200 0.6525 0.5775 0.7725 ;
        VIA 0.8925 0.3375 VIA12_slot ;
        VIA 0.8925 0.7125 VIA12_slot ;
        VIA 0.5775 0.3375 VIA12_slot ;
        VIA 0.5775 0.7125 VIA12_slot ;
        END
    END ZN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1425 0.4725 1.3350 0.5475 ;
        RECT 0.0675 0.3675 0.1425 0.6825 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.4250 -0.0750 1.4700 0.0750 ;
        RECT 1.3050 -0.0750 1.4250 0.2925 ;
        RECT 1.0050 -0.0750 1.3050 0.0750 ;
        RECT 0.8850 -0.0750 1.0050 0.2025 ;
        RECT 0.5850 -0.0750 0.8850 0.0750 ;
        RECT 0.4650 -0.0750 0.5850 0.2025 ;
        RECT 0.1425 -0.0750 0.4650 0.0750 ;
        RECT 0.0675 -0.0750 0.1425 0.2475 ;
        RECT 0.0000 -0.0750 0.0675 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.4250 0.9750 1.4700 1.1250 ;
        RECT 1.3050 0.6600 1.4250 1.1250 ;
        RECT 1.0050 0.9750 1.3050 1.1250 ;
        RECT 0.8850 0.8475 1.0050 1.1250 ;
        RECT 0.5850 0.9750 0.8850 1.1250 ;
        RECT 0.4650 0.8475 0.5850 1.1250 ;
        RECT 0.1425 0.9750 0.4650 1.1250 ;
        RECT 0.0675 0.8025 0.1425 1.1250 ;
        RECT 0.0000 0.9750 0.0675 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.3350 0.2250 1.3950 0.2850 ;
        RECT 1.3350 0.6675 1.3950 0.7275 ;
        RECT 1.3350 0.8325 1.3950 0.8925 ;
        RECT 1.2300 0.4800 1.2900 0.5400 ;
        RECT 1.1250 0.3075 1.1850 0.3675 ;
        RECT 1.1250 0.6825 1.1850 0.7425 ;
        RECT 1.0200 0.4800 1.0800 0.5400 ;
        RECT 0.9150 0.1350 0.9750 0.1950 ;
        RECT 0.9150 0.8550 0.9750 0.9150 ;
        RECT 0.8100 0.4800 0.8700 0.5400 ;
        RECT 0.7050 0.3075 0.7650 0.3675 ;
        RECT 0.7050 0.6825 0.7650 0.7425 ;
        RECT 0.6000 0.4800 0.6600 0.5400 ;
        RECT 0.4950 0.1350 0.5550 0.1950 ;
        RECT 0.4950 0.8550 0.5550 0.9150 ;
        RECT 0.3900 0.4800 0.4500 0.5400 ;
        RECT 0.2850 0.3075 0.3450 0.3675 ;
        RECT 0.2850 0.6825 0.3450 0.7425 ;
        RECT 0.1800 0.4800 0.2400 0.5400 ;
        RECT 0.0750 0.1575 0.1350 0.2175 ;
        RECT 0.0750 0.8325 0.1350 0.8925 ;
        LAYER M1 ;
        RECT 0.2775 0.2775 1.2000 0.3975 ;
        RECT 0.2775 0.6525 1.2000 0.7725 ;
        LAYER M2 ;
        RECT 0.9225 0.2775 1.0500 0.3975 ;
        RECT 0.9225 0.6525 1.0500 0.7725 ;
        RECT 0.4200 0.2775 0.5475 0.3975 ;
        RECT 0.4200 0.6525 0.5475 0.7725 ;
    END
END INV_0110


MACRO INV_0111
    CLASS CORE ;
    FOREIGN INV_0111 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.0500 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 0.3675 0.2700 0.6825 0.7800 ;
        VIA 0.5250 0.3525 VIA12_slot ;
        VIA 0.5250 0.6975 VIA12_slot ;
        END
    END ZN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1425 0.4725 0.9150 0.5475 ;
        RECT 0.0675 0.3675 0.1425 0.6825 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.0050 -0.0750 1.0500 0.0750 ;
        RECT 0.8850 -0.0750 1.0050 0.2925 ;
        RECT 0.5850 -0.0750 0.8850 0.0750 ;
        RECT 0.4650 -0.0750 0.5850 0.2025 ;
        RECT 0.1425 -0.0750 0.4650 0.0750 ;
        RECT 0.0675 -0.0750 0.1425 0.2475 ;
        RECT 0.0000 -0.0750 0.0675 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.0050 0.9750 1.0500 1.1250 ;
        RECT 0.8850 0.6600 1.0050 1.1250 ;
        RECT 0.5850 0.9750 0.8850 1.1250 ;
        RECT 0.4650 0.8475 0.5850 1.1250 ;
        RECT 0.1425 0.9750 0.4650 1.1250 ;
        RECT 0.0675 0.8025 0.1425 1.1250 ;
        RECT 0.0000 0.9750 0.0675 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 0.9150 0.2175 0.9750 0.2775 ;
        RECT 0.9150 0.6675 0.9750 0.7275 ;
        RECT 0.9150 0.8325 0.9750 0.8925 ;
        RECT 0.8100 0.4800 0.8700 0.5400 ;
        RECT 0.7050 0.3075 0.7650 0.3675 ;
        RECT 0.7050 0.6825 0.7650 0.7425 ;
        RECT 0.6000 0.4800 0.6600 0.5400 ;
        RECT 0.4950 0.1350 0.5550 0.1950 ;
        RECT 0.4950 0.8550 0.5550 0.9150 ;
        RECT 0.3900 0.4800 0.4500 0.5400 ;
        RECT 0.2850 0.3075 0.3450 0.3675 ;
        RECT 0.2850 0.6825 0.3450 0.7425 ;
        RECT 0.1800 0.4800 0.2400 0.5400 ;
        RECT 0.0750 0.1575 0.1350 0.2175 ;
        RECT 0.0750 0.8325 0.1350 0.8925 ;
        LAYER M1 ;
        RECT 0.2775 0.2775 0.7800 0.3975 ;
        RECT 0.2775 0.6525 0.7800 0.7725 ;
    END
END INV_0111


MACRO INV_1000
    CLASS CORE ;
    FOREIGN INV_1000 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.4200 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.3075 0.1500 0.3825 0.9000 ;
        RECT 0.2550 0.1500 0.3075 0.2550 ;
        RECT 0.2625 0.6675 0.3075 0.9000 ;
        END
    END ZN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1425 0.4425 0.2325 0.5925 ;
        RECT 0.0675 0.3675 0.1425 0.6825 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.1650 -0.0750 0.4200 0.0750 ;
        RECT 0.0450 -0.0750 0.1650 0.2325 ;
        RECT 0.0000 -0.0750 0.0450 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.1650 0.9750 0.4200 1.1250 ;
        RECT 0.0450 0.8175 0.1650 1.1250 ;
        RECT 0.0000 0.9750 0.0450 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 0.2850 0.1575 0.3450 0.2175 ;
        RECT 0.2850 0.8175 0.3450 0.8775 ;
        RECT 0.1725 0.4875 0.2325 0.5475 ;
        RECT 0.0750 0.1575 0.1350 0.2175 ;
        RECT 0.0750 0.8325 0.1350 0.8925 ;
    END
END INV_1000


MACRO INV_1010
    CLASS CORE ;
    FOREIGN INV_1010 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.4200 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.3075 0.2025 0.3825 0.8475 ;
        RECT 0.2775 0.2025 0.3075 0.3825 ;
        RECT 0.2775 0.6675 0.3075 0.8475 ;
        END
    END ZN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1425 0.4425 0.2325 0.5925 ;
        RECT 0.0675 0.3675 0.1425 0.6825 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.1425 -0.0750 0.4200 0.0750 ;
        RECT 0.0675 -0.0750 0.1425 0.2475 ;
        RECT 0.0000 -0.0750 0.0675 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.1425 0.9750 0.4200 1.1250 ;
        RECT 0.0675 0.8025 0.1425 1.1250 ;
        RECT 0.0000 0.9750 0.0675 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 0.2850 0.2475 0.3450 0.3075 ;
        RECT 0.2850 0.7425 0.3450 0.8025 ;
        RECT 0.1725 0.4875 0.2325 0.5475 ;
        RECT 0.0750 0.1575 0.1350 0.2175 ;
        RECT 0.0750 0.8325 0.1350 0.8925 ;
    END
END INV_1010


MACRO INV_1100
    CLASS CORE ;
    FOREIGN INV_1100 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.5700 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 1.9425 0.2775 2.1000 0.3975 ;
        RECT 1.9425 0.6525 2.1000 0.7725 ;
        RECT 1.6275 0.2775 1.9425 0.7725 ;
        RECT 1.4700 0.2775 1.6275 0.3975 ;
        RECT 1.4700 0.6525 1.6275 0.7725 ;
        VIA 1.9425 0.3375 VIA12_slot ;
        VIA 1.9425 0.7125 VIA12_slot ;
        VIA 1.6275 0.3375 VIA12_slot ;
        VIA 1.6275 0.7125 VIA12_slot ;
        END
    END ZN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1425 0.4725 3.4650 0.5475 ;
        RECT 0.0675 0.3675 0.1425 0.6825 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 3.5250 -0.0750 3.5700 0.0750 ;
        RECT 3.4050 -0.0750 3.5250 0.2925 ;
        RECT 3.1050 -0.0750 3.4050 0.0750 ;
        RECT 2.9850 -0.0750 3.1050 0.2025 ;
        RECT 2.6850 -0.0750 2.9850 0.0750 ;
        RECT 2.5650 -0.0750 2.6850 0.2025 ;
        RECT 2.2650 -0.0750 2.5650 0.0750 ;
        RECT 2.1450 -0.0750 2.2650 0.2025 ;
        RECT 1.8450 -0.0750 2.1450 0.0750 ;
        RECT 1.7250 -0.0750 1.8450 0.2025 ;
        RECT 1.4250 -0.0750 1.7250 0.0750 ;
        RECT 1.3050 -0.0750 1.4250 0.2025 ;
        RECT 1.0050 -0.0750 1.3050 0.0750 ;
        RECT 0.8850 -0.0750 1.0050 0.2025 ;
        RECT 0.5850 -0.0750 0.8850 0.0750 ;
        RECT 0.4650 -0.0750 0.5850 0.2025 ;
        RECT 0.1425 -0.0750 0.4650 0.0750 ;
        RECT 0.0675 -0.0750 0.1425 0.2475 ;
        RECT 0.0000 -0.0750 0.0675 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 3.5250 0.9750 3.5700 1.1250 ;
        RECT 3.4050 0.6600 3.5250 1.1250 ;
        RECT 3.1050 0.9750 3.4050 1.1250 ;
        RECT 2.9850 0.8475 3.1050 1.1250 ;
        RECT 2.6850 0.9750 2.9850 1.1250 ;
        RECT 2.5650 0.8475 2.6850 1.1250 ;
        RECT 2.2650 0.9750 2.5650 1.1250 ;
        RECT 2.1450 0.8475 2.2650 1.1250 ;
        RECT 1.8450 0.9750 2.1450 1.1250 ;
        RECT 1.7250 0.8475 1.8450 1.1250 ;
        RECT 1.4250 0.9750 1.7250 1.1250 ;
        RECT 1.3050 0.8475 1.4250 1.1250 ;
        RECT 1.0050 0.9750 1.3050 1.1250 ;
        RECT 0.8850 0.8475 1.0050 1.1250 ;
        RECT 0.5850 0.9750 0.8850 1.1250 ;
        RECT 0.4650 0.8475 0.5850 1.1250 ;
        RECT 0.1425 0.9750 0.4650 1.1250 ;
        RECT 0.0675 0.8025 0.1425 1.1250 ;
        RECT 0.0000 0.9750 0.0675 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 3.4350 0.2175 3.4950 0.2775 ;
        RECT 3.4350 0.6675 3.4950 0.7275 ;
        RECT 3.4350 0.8325 3.4950 0.8925 ;
        RECT 3.3300 0.4800 3.3900 0.5400 ;
        RECT 3.2250 0.3075 3.2850 0.3675 ;
        RECT 3.2250 0.6825 3.2850 0.7425 ;
        RECT 3.1200 0.4800 3.1800 0.5400 ;
        RECT 3.0150 0.1350 3.0750 0.1950 ;
        RECT 3.0150 0.8550 3.0750 0.9150 ;
        RECT 2.9100 0.4800 2.9700 0.5400 ;
        RECT 2.8050 0.3075 2.8650 0.3675 ;
        RECT 2.8050 0.6825 2.8650 0.7425 ;
        RECT 2.7000 0.4800 2.7600 0.5400 ;
        RECT 2.5950 0.1350 2.6550 0.1950 ;
        RECT 2.5950 0.8550 2.6550 0.9150 ;
        RECT 2.4900 0.4800 2.5500 0.5400 ;
        RECT 2.3850 0.3075 2.4450 0.3675 ;
        RECT 2.3850 0.6825 2.4450 0.7425 ;
        RECT 2.2800 0.4800 2.3400 0.5400 ;
        RECT 2.1750 0.1350 2.2350 0.1950 ;
        RECT 2.1750 0.8550 2.2350 0.9150 ;
        RECT 2.0700 0.4800 2.1300 0.5400 ;
        RECT 1.9650 0.3075 2.0250 0.3675 ;
        RECT 1.9650 0.6825 2.0250 0.7425 ;
        RECT 1.8600 0.4800 1.9200 0.5400 ;
        RECT 1.7550 0.1350 1.8150 0.1950 ;
        RECT 1.7550 0.8550 1.8150 0.9150 ;
        RECT 1.6500 0.4800 1.7100 0.5400 ;
        RECT 1.5450 0.3075 1.6050 0.3675 ;
        RECT 1.5450 0.6825 1.6050 0.7425 ;
        RECT 1.4400 0.4800 1.5000 0.5400 ;
        RECT 1.3350 0.1350 1.3950 0.1950 ;
        RECT 1.3350 0.8550 1.3950 0.9150 ;
        RECT 1.2300 0.4800 1.2900 0.5400 ;
        RECT 1.1250 0.3075 1.1850 0.3675 ;
        RECT 1.1250 0.6825 1.1850 0.7425 ;
        RECT 1.0200 0.4800 1.0800 0.5400 ;
        RECT 0.9150 0.1350 0.9750 0.1950 ;
        RECT 0.9150 0.8550 0.9750 0.9150 ;
        RECT 0.8100 0.4800 0.8700 0.5400 ;
        RECT 0.7050 0.3075 0.7650 0.3675 ;
        RECT 0.7050 0.6825 0.7650 0.7425 ;
        RECT 0.6000 0.4800 0.6600 0.5400 ;
        RECT 0.4950 0.1350 0.5550 0.1950 ;
        RECT 0.4950 0.8550 0.5550 0.9150 ;
        RECT 0.3900 0.4800 0.4500 0.5400 ;
        RECT 0.2850 0.3075 0.3450 0.3675 ;
        RECT 0.2850 0.6825 0.3450 0.7425 ;
        RECT 0.1800 0.4800 0.2400 0.5400 ;
        RECT 0.0750 0.1575 0.1350 0.2175 ;
        RECT 0.0750 0.8325 0.1350 0.8925 ;
        LAYER M1 ;
        RECT 0.2775 0.2775 3.3000 0.3975 ;
        RECT 0.2775 0.6525 3.3000 0.7725 ;
        LAYER M2 ;
        RECT 1.9725 0.2775 2.1000 0.3975 ;
        RECT 1.9725 0.6525 2.1000 0.7725 ;
        RECT 1.4700 0.2775 1.5975 0.3975 ;
        RECT 1.4700 0.6525 1.5975 0.7725 ;
    END
END INV_1100


MACRO LHQ_0011
    CLASS CORE ;
    FOREIGN LHQ_0011 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.3100 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 2.1975 0.3075 2.2725 0.7425 ;
        RECT 2.0325 0.3075 2.1975 0.3825 ;
        RECT 2.0325 0.6675 2.1975 0.7425 ;
        RECT 1.9575 0.2100 2.0325 0.3825 ;
        RECT 1.9575 0.6675 2.0325 0.8475 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.4575 0.8625 0.6675 0.9375 ;
        RECT 0.3525 0.5700 0.4575 0.9375 ;
        RECT 0.1050 0.8625 0.3525 0.9375 ;
        VIA 0.4050 0.6450 VIA12_square ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.6275 0.1125 1.7400 0.4125 ;
        RECT 1.1625 0.1125 1.6275 0.1875 ;
        VIA 1.6875 0.3375 VIA12_square ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 2.2650 -0.0750 2.3100 0.0750 ;
        RECT 2.1450 -0.0750 2.2650 0.2325 ;
        RECT 1.8450 -0.0750 2.1450 0.0750 ;
        RECT 1.7250 -0.0750 1.8450 0.1800 ;
        RECT 1.0050 -0.0750 1.7250 0.0750 ;
        RECT 0.8850 -0.0750 1.0050 0.1800 ;
        RECT 0.3750 -0.0750 0.8850 0.0750 ;
        RECT 0.2550 -0.0750 0.3750 0.1875 ;
        RECT 0.0000 -0.0750 0.2550 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 2.2650 0.9750 2.3100 1.1250 ;
        RECT 2.1450 0.8175 2.2650 1.1250 ;
        RECT 1.8600 0.9750 2.1450 1.1250 ;
        RECT 1.7550 0.8400 1.8600 1.1250 ;
        RECT 1.0050 0.9750 1.7550 1.1250 ;
        RECT 0.8850 0.8700 1.0050 1.1250 ;
        RECT 0.3600 0.9750 0.8850 1.1250 ;
        RECT 0.2550 0.8100 0.3600 1.1250 ;
        RECT 0.0000 0.9750 0.2550 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 2.1750 0.1575 2.2350 0.2175 ;
        RECT 2.1750 0.8325 2.2350 0.8925 ;
        RECT 2.0625 0.4950 2.1225 0.5550 ;
        RECT 1.9650 0.2400 2.0250 0.3000 ;
        RECT 1.9650 0.7575 2.0250 0.8175 ;
        RECT 1.8600 0.4875 1.9200 0.5475 ;
        RECT 1.7550 0.1200 1.8150 0.1800 ;
        RECT 1.7550 0.8700 1.8150 0.9300 ;
        RECT 1.6425 0.4425 1.7025 0.5025 ;
        RECT 1.4475 0.4200 1.5075 0.4800 ;
        RECT 1.4400 0.6600 1.5000 0.7200 ;
        RECT 1.3350 0.1575 1.3950 0.2175 ;
        RECT 1.3350 0.8325 1.3950 0.8925 ;
        RECT 1.2225 0.3300 1.2825 0.3900 ;
        RECT 1.2225 0.6600 1.2825 0.7200 ;
        RECT 1.0125 0.4875 1.0725 0.5475 ;
        RECT 0.9150 0.1200 0.9750 0.1800 ;
        RECT 0.9150 0.8700 0.9750 0.9300 ;
        RECT 0.8025 0.4950 0.8625 0.5550 ;
        RECT 0.7050 0.2325 0.7650 0.2925 ;
        RECT 0.7050 0.7500 0.7650 0.8100 ;
        RECT 0.4950 0.1800 0.5550 0.2400 ;
        RECT 0.4950 0.8325 0.5550 0.8925 ;
        RECT 0.3825 0.3975 0.4425 0.4575 ;
        RECT 0.2850 0.1275 0.3450 0.1875 ;
        RECT 0.2850 0.8400 0.3450 0.9000 ;
        RECT 0.1875 0.5925 0.2475 0.6525 ;
        RECT 0.0750 0.1725 0.1350 0.2325 ;
        RECT 0.0750 0.8100 0.1350 0.8700 ;
        LAYER M1 ;
        RECT 1.8825 0.4650 2.1225 0.5850 ;
        RECT 1.8075 0.4650 1.8825 0.6825 ;
        RECT 1.7325 0.2550 1.8600 0.3675 ;
        RECT 1.6275 0.2550 1.7325 0.5400 ;
        RECT 1.4625 0.6300 1.6800 0.7200 ;
        RECT 1.5300 0.7950 1.6800 0.9000 ;
        RECT 1.3875 0.1500 1.5525 0.3450 ;
        RECT 1.4175 0.4200 1.5375 0.5550 ;
        RECT 1.2900 0.8250 1.5300 0.9000 ;
        RECT 1.3575 0.6300 1.4625 0.7500 ;
        RECT 1.2825 0.4800 1.4175 0.5550 ;
        RECT 1.2975 0.1500 1.3875 0.2250 ;
        RECT 1.1925 0.3000 1.3125 0.4050 ;
        RECT 1.2075 0.4800 1.2825 0.7500 ;
        RECT 1.1625 0.6300 1.2075 0.7500 ;
        RECT 1.0875 0.1500 1.1925 0.4050 ;
        RECT 1.0875 0.6300 1.1625 0.8325 ;
        RECT 1.0125 0.4800 1.1025 0.5550 ;
        RECT 0.9375 0.2625 1.0125 0.7950 ;
        RECT 0.7950 0.2625 0.9375 0.3375 ;
        RECT 0.7725 0.7200 0.9375 0.7950 ;
        RECT 0.6675 0.4125 0.8625 0.6450 ;
        RECT 0.7050 0.1950 0.7950 0.3375 ;
        RECT 0.6975 0.7200 0.7725 0.8700 ;
        RECT 0.5175 0.1500 0.5925 0.9000 ;
        RECT 0.4875 0.1500 0.5175 0.2700 ;
        RECT 0.4650 0.8100 0.5175 0.9000 ;
        RECT 0.4125 0.3675 0.4425 0.4875 ;
        RECT 0.3375 0.5625 0.4425 0.7350 ;
        RECT 0.3375 0.2625 0.4125 0.4875 ;
        RECT 0.1575 0.2625 0.3375 0.3375 ;
        RECT 0.1875 0.5625 0.3375 0.6825 ;
        RECT 0.1125 0.1500 0.1575 0.3375 ;
        RECT 0.1125 0.7800 0.1575 0.9000 ;
        RECT 0.0375 0.1500 0.1125 0.9000 ;
        LAYER VIA1 ;
        RECT 1.8075 0.5625 1.8825 0.6375 ;
        RECT 1.5675 0.8100 1.6425 0.8850 ;
        RECT 1.4325 0.2625 1.5075 0.3375 ;
        RECT 1.4025 0.6450 1.4775 0.7200 ;
        RECT 1.1025 0.2625 1.1775 0.3375 ;
        RECT 1.0875 0.6750 1.1625 0.7500 ;
        RECT 0.7275 0.5625 0.8025 0.6375 ;
        RECT 0.5175 0.4125 0.5925 0.4875 ;
        RECT 0.2925 0.2625 0.3675 0.3375 ;
        LAYER M2 ;
        RECT 1.7475 0.5625 1.9650 0.6375 ;
        RECT 1.6725 0.4950 1.7475 0.8850 ;
        RECT 1.5525 0.4950 1.6725 0.5700 ;
        RECT 1.5750 0.8100 1.6725 0.8850 ;
        RECT 1.4775 0.8100 1.5750 0.9375 ;
        RECT 1.4775 0.2625 1.5525 0.5700 ;
        RECT 1.3275 0.6450 1.5525 0.7200 ;
        RECT 1.3425 0.2625 1.4775 0.3375 ;
        RECT 0.8625 0.8625 1.4775 0.9375 ;
        RECT 1.2525 0.4125 1.3275 0.7200 ;
        RECT 1.2225 0.4125 1.2525 0.4875 ;
        RECT 1.1475 0.2625 1.2225 0.4875 ;
        RECT 1.0125 0.6375 1.1775 0.7875 ;
        RECT 0.2475 0.2625 1.1475 0.3375 ;
        RECT 0.9375 0.4125 1.0125 0.7875 ;
        RECT 0.4425 0.4125 0.9375 0.4875 ;
        RECT 0.7875 0.5625 0.8625 0.9375 ;
        RECT 0.6525 0.5625 0.7875 0.6375 ;
    END
END LHQ_0011


MACRO LHQ_0111
    CLASS CORE ;
    FOREIGN LHQ_0111 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.7300 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 2.0475 0.2325 2.3625 0.7350 ;
        VIA 2.2050 0.3150 VIA12_slot ;
        VIA 2.2050 0.6525 VIA12_slot ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.4575 0.8625 0.6675 0.9375 ;
        RECT 0.3525 0.5700 0.4575 0.9375 ;
        RECT 0.1050 0.8625 0.3525 0.9375 ;
        VIA 0.4050 0.6450 VIA12_square ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.6275 0.1125 1.7400 0.4125 ;
        RECT 1.1625 0.1125 1.6275 0.1875 ;
        VIA 1.6875 0.3375 VIA12_square ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 2.6625 -0.0750 2.7300 0.0750 ;
        RECT 2.5875 -0.0750 2.6625 0.2475 ;
        RECT 2.2650 -0.0750 2.5875 0.0750 ;
        RECT 2.1450 -0.0750 2.2650 0.1875 ;
        RECT 1.8450 -0.0750 2.1450 0.0750 ;
        RECT 1.7250 -0.0750 1.8450 0.1800 ;
        RECT 1.0050 -0.0750 1.7250 0.0750 ;
        RECT 0.8850 -0.0750 1.0050 0.1800 ;
        RECT 0.3750 -0.0750 0.8850 0.0750 ;
        RECT 0.2550 -0.0750 0.3750 0.1875 ;
        RECT 0.0000 -0.0750 0.2550 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 2.6850 0.9750 2.7300 1.1250 ;
        RECT 2.5650 0.6450 2.6850 1.1250 ;
        RECT 2.2650 0.9750 2.5650 1.1250 ;
        RECT 2.1450 0.8175 2.2650 1.1250 ;
        RECT 1.8600 0.9750 2.1450 1.1250 ;
        RECT 1.7550 0.8400 1.8600 1.1250 ;
        RECT 1.0050 0.9750 1.7550 1.1250 ;
        RECT 0.8850 0.8700 1.0050 1.1250 ;
        RECT 0.3600 0.9750 0.8850 1.1250 ;
        RECT 0.2550 0.8100 0.3600 1.1250 ;
        RECT 0.0000 0.9750 0.2550 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 2.5950 0.1575 2.6550 0.2175 ;
        RECT 2.5950 0.6675 2.6550 0.7275 ;
        RECT 2.5950 0.8325 2.6550 0.8925 ;
        RECT 2.4900 0.4725 2.5500 0.5325 ;
        RECT 2.3850 0.2850 2.4450 0.3450 ;
        RECT 2.3850 0.6525 2.4450 0.7125 ;
        RECT 2.2800 0.4725 2.3400 0.5325 ;
        RECT 2.1750 0.1275 2.2350 0.1875 ;
        RECT 2.1750 0.8325 2.2350 0.8925 ;
        RECT 2.0700 0.4725 2.1300 0.5325 ;
        RECT 1.9650 0.2700 2.0250 0.3300 ;
        RECT 1.9650 0.6525 2.0250 0.7125 ;
        RECT 1.8600 0.4725 1.9200 0.5325 ;
        RECT 1.7550 0.1200 1.8150 0.1800 ;
        RECT 1.7550 0.8700 1.8150 0.9300 ;
        RECT 1.6425 0.4425 1.7025 0.5025 ;
        RECT 1.4475 0.4200 1.5075 0.4800 ;
        RECT 1.4400 0.6600 1.5000 0.7200 ;
        RECT 1.3350 0.1575 1.3950 0.2175 ;
        RECT 1.3350 0.8325 1.3950 0.8925 ;
        RECT 1.2225 0.3300 1.2825 0.3900 ;
        RECT 1.2225 0.6600 1.2825 0.7200 ;
        RECT 1.0125 0.4875 1.0725 0.5475 ;
        RECT 0.9150 0.1200 0.9750 0.1800 ;
        RECT 0.9150 0.8700 0.9750 0.9300 ;
        RECT 0.8025 0.4950 0.8625 0.5550 ;
        RECT 0.7050 0.2325 0.7650 0.2925 ;
        RECT 0.7050 0.7500 0.7650 0.8100 ;
        RECT 0.4950 0.1800 0.5550 0.2400 ;
        RECT 0.4950 0.8325 0.5550 0.8925 ;
        RECT 0.3825 0.3975 0.4425 0.4575 ;
        RECT 0.2850 0.1275 0.3450 0.1875 ;
        RECT 0.2850 0.8400 0.3450 0.9000 ;
        RECT 0.1875 0.5925 0.2475 0.6525 ;
        RECT 0.0750 0.1725 0.1350 0.2325 ;
        RECT 0.0750 0.8100 0.1350 0.8700 ;
        LAYER M1 ;
        RECT 1.8825 0.4650 2.5800 0.5400 ;
        RECT 2.0475 0.2625 2.4750 0.3600 ;
        RECT 1.9650 0.6150 2.4675 0.7425 ;
        RECT 1.9650 0.2400 2.0475 0.3600 ;
        RECT 1.8075 0.4650 1.8825 0.6825 ;
        RECT 1.7325 0.2550 1.8600 0.3675 ;
        RECT 1.6275 0.2550 1.7325 0.5400 ;
        RECT 1.4625 0.6300 1.6800 0.7200 ;
        RECT 1.5300 0.7950 1.6800 0.9000 ;
        RECT 1.3875 0.1500 1.5525 0.3450 ;
        RECT 1.4175 0.4200 1.5375 0.5550 ;
        RECT 1.2900 0.8250 1.5300 0.9000 ;
        RECT 1.3575 0.6300 1.4625 0.7500 ;
        RECT 1.2825 0.4800 1.4175 0.5550 ;
        RECT 1.2975 0.1500 1.3875 0.2250 ;
        RECT 1.1925 0.3000 1.3125 0.4050 ;
        RECT 1.2075 0.4800 1.2825 0.7500 ;
        RECT 1.1625 0.6300 1.2075 0.7500 ;
        RECT 1.0875 0.1500 1.1925 0.4050 ;
        RECT 1.0875 0.6300 1.1625 0.8325 ;
        RECT 1.0125 0.4800 1.1025 0.5550 ;
        RECT 0.9375 0.2625 1.0125 0.7950 ;
        RECT 0.7950 0.2625 0.9375 0.3375 ;
        RECT 0.7725 0.7200 0.9375 0.7950 ;
        RECT 0.6675 0.4125 0.8625 0.6450 ;
        RECT 0.7050 0.1950 0.7950 0.3375 ;
        RECT 0.6975 0.7200 0.7725 0.8700 ;
        RECT 0.5175 0.1500 0.5925 0.9000 ;
        RECT 0.4875 0.1500 0.5175 0.2700 ;
        RECT 0.4650 0.8100 0.5175 0.9000 ;
        RECT 0.4125 0.3675 0.4425 0.4875 ;
        RECT 0.3375 0.5625 0.4425 0.7350 ;
        RECT 0.3375 0.2625 0.4125 0.4875 ;
        RECT 0.1575 0.2625 0.3375 0.3375 ;
        RECT 0.1875 0.5625 0.3375 0.6825 ;
        RECT 0.1125 0.1500 0.1575 0.3375 ;
        RECT 0.1125 0.7800 0.1575 0.9000 ;
        RECT 0.0375 0.1500 0.1125 0.9000 ;
        LAYER VIA1 ;
        RECT 1.8075 0.5625 1.8825 0.6375 ;
        RECT 1.5675 0.8100 1.6425 0.8850 ;
        RECT 1.4325 0.2625 1.5075 0.3375 ;
        RECT 1.4025 0.6450 1.4775 0.7200 ;
        RECT 1.1025 0.2625 1.1775 0.3375 ;
        RECT 1.0875 0.6750 1.1625 0.7500 ;
        RECT 0.7275 0.5625 0.8025 0.6375 ;
        RECT 0.5175 0.4125 0.5925 0.4875 ;
        RECT 0.2925 0.2625 0.3675 0.3375 ;
        LAYER M2 ;
        RECT 1.8075 0.4950 1.8825 0.8850 ;
        RECT 1.5525 0.4950 1.8075 0.5700 ;
        RECT 1.5750 0.8100 1.8075 0.8850 ;
        RECT 1.4775 0.8100 1.5750 0.9375 ;
        RECT 1.4775 0.2625 1.5525 0.5700 ;
        RECT 1.3275 0.6450 1.5525 0.7200 ;
        RECT 1.3425 0.2625 1.4775 0.3375 ;
        RECT 0.8625 0.8625 1.4775 0.9375 ;
        RECT 1.2525 0.4125 1.3275 0.7200 ;
        RECT 1.2225 0.4125 1.2525 0.4875 ;
        RECT 1.1475 0.2625 1.2225 0.4875 ;
        RECT 1.0125 0.6375 1.1775 0.7875 ;
        RECT 0.2475 0.2625 1.1475 0.3375 ;
        RECT 0.9375 0.4125 1.0125 0.7875 ;
        RECT 0.4425 0.4125 0.9375 0.4875 ;
        RECT 0.7875 0.5625 0.8625 0.9375 ;
        RECT 0.6525 0.5625 0.7875 0.6375 ;
    END
END LHQ_0111


MACRO LHQ_1010
    CLASS CORE ;
    FOREIGN LHQ_1010 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.1000 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 1.9875 0.2175 2.0625 0.8325 ;
        RECT 1.9575 0.2175 1.9875 0.3825 ;
        RECT 1.9650 0.6675 1.9875 0.8325 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.4575 0.8625 0.6675 0.9375 ;
        RECT 0.3525 0.5700 0.4575 0.9375 ;
        RECT 0.1050 0.8625 0.3525 0.9375 ;
        VIA 0.4050 0.6450 VIA12_square ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.6275 0.1125 1.7400 0.4125 ;
        RECT 1.1625 0.1125 1.6275 0.1875 ;
        VIA 1.6875 0.3375 VIA12_square ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.8450 -0.0750 2.1000 0.0750 ;
        RECT 1.7250 -0.0750 1.8450 0.1800 ;
        RECT 1.0050 -0.0750 1.7250 0.0750 ;
        RECT 0.8850 -0.0750 1.0050 0.1800 ;
        RECT 0.3750 -0.0750 0.8850 0.0750 ;
        RECT 0.2550 -0.0750 0.3750 0.1875 ;
        RECT 0.0000 -0.0750 0.2550 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.8600 0.9750 2.1000 1.1250 ;
        RECT 1.7550 0.8400 1.8600 1.1250 ;
        RECT 1.0050 0.9750 1.7550 1.1250 ;
        RECT 0.8850 0.8700 1.0050 1.1250 ;
        RECT 0.3600 0.9750 0.8850 1.1250 ;
        RECT 0.2550 0.8100 0.3600 1.1250 ;
        RECT 0.0000 0.9750 0.2550 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.9650 0.2700 2.0250 0.3300 ;
        RECT 1.9650 0.7200 2.0250 0.7800 ;
        RECT 1.8525 0.4725 1.9125 0.5325 ;
        RECT 1.7550 0.1200 1.8150 0.1800 ;
        RECT 1.7550 0.8700 1.8150 0.9300 ;
        RECT 1.6425 0.4425 1.7025 0.5025 ;
        RECT 1.4475 0.4200 1.5075 0.4800 ;
        RECT 1.4400 0.6600 1.5000 0.7200 ;
        RECT 1.3350 0.1575 1.3950 0.2175 ;
        RECT 1.3350 0.8325 1.3950 0.8925 ;
        RECT 1.2225 0.3300 1.2825 0.3900 ;
        RECT 1.2225 0.6600 1.2825 0.7200 ;
        RECT 1.0125 0.4875 1.0725 0.5475 ;
        RECT 0.9150 0.1200 0.9750 0.1800 ;
        RECT 0.9150 0.8700 0.9750 0.9300 ;
        RECT 0.8025 0.4950 0.8625 0.5550 ;
        RECT 0.7050 0.2325 0.7650 0.2925 ;
        RECT 0.7050 0.7500 0.7650 0.8100 ;
        RECT 0.4950 0.1800 0.5550 0.2400 ;
        RECT 0.4950 0.8325 0.5550 0.8925 ;
        RECT 0.3825 0.3975 0.4425 0.4575 ;
        RECT 0.2850 0.1275 0.3450 0.1875 ;
        RECT 0.2850 0.8400 0.3450 0.9000 ;
        RECT 0.1875 0.5925 0.2475 0.6525 ;
        RECT 0.0750 0.1725 0.1350 0.2325 ;
        RECT 0.0750 0.8100 0.1350 0.8700 ;
        LAYER M1 ;
        RECT 1.8900 0.4425 1.9125 0.6075 ;
        RECT 1.8075 0.4425 1.8900 0.7650 ;
        RECT 1.7325 0.2550 1.8600 0.3675 ;
        RECT 1.7850 0.6000 1.8075 0.7650 ;
        RECT 1.6275 0.2550 1.7325 0.5400 ;
        RECT 1.4625 0.6300 1.6800 0.7200 ;
        RECT 1.5300 0.7950 1.6800 0.9000 ;
        RECT 1.3875 0.1500 1.5525 0.3450 ;
        RECT 1.4175 0.4200 1.5375 0.5550 ;
        RECT 1.2900 0.8250 1.5300 0.9000 ;
        RECT 1.3575 0.6300 1.4625 0.7500 ;
        RECT 1.2825 0.4800 1.4175 0.5550 ;
        RECT 1.2975 0.1500 1.3875 0.2250 ;
        RECT 1.1925 0.3000 1.3125 0.4050 ;
        RECT 1.2075 0.4800 1.2825 0.7500 ;
        RECT 1.1625 0.6300 1.2075 0.7500 ;
        RECT 1.0875 0.1500 1.1925 0.4050 ;
        RECT 1.0875 0.6300 1.1625 0.8325 ;
        RECT 1.0125 0.4800 1.1025 0.5550 ;
        RECT 0.9375 0.2625 1.0125 0.7950 ;
        RECT 0.7950 0.2625 0.9375 0.3375 ;
        RECT 0.7725 0.7200 0.9375 0.7950 ;
        RECT 0.6675 0.4125 0.8625 0.6450 ;
        RECT 0.7050 0.1950 0.7950 0.3375 ;
        RECT 0.6975 0.7200 0.7725 0.8700 ;
        RECT 0.5175 0.1500 0.5925 0.9000 ;
        RECT 0.4875 0.1500 0.5175 0.2700 ;
        RECT 0.4650 0.8100 0.5175 0.9000 ;
        RECT 0.4125 0.3675 0.4425 0.4875 ;
        RECT 0.3375 0.5625 0.4425 0.7350 ;
        RECT 0.3375 0.2625 0.4125 0.4875 ;
        RECT 0.1575 0.2625 0.3375 0.3375 ;
        RECT 0.1875 0.5625 0.3375 0.6825 ;
        RECT 0.1125 0.1500 0.1575 0.3375 ;
        RECT 0.1125 0.7800 0.1575 0.9000 ;
        RECT 0.0375 0.1500 0.1125 0.9000 ;
        LAYER VIA1 ;
        RECT 1.8150 0.5625 1.8900 0.6375 ;
        RECT 1.5675 0.8100 1.6425 0.8850 ;
        RECT 1.4325 0.2625 1.5075 0.3375 ;
        RECT 1.4025 0.6450 1.4775 0.7200 ;
        RECT 1.1025 0.2625 1.1775 0.3375 ;
        RECT 1.0875 0.6750 1.1625 0.7500 ;
        RECT 0.7275 0.5625 0.8025 0.6375 ;
        RECT 0.5175 0.4125 0.5925 0.4875 ;
        RECT 0.2925 0.2625 0.3675 0.3375 ;
        LAYER M2 ;
        RECT 1.7475 0.5625 1.9650 0.6375 ;
        RECT 1.6725 0.4950 1.7475 0.8850 ;
        RECT 1.5525 0.4950 1.6725 0.5700 ;
        RECT 1.5750 0.8100 1.6725 0.8850 ;
        RECT 1.4775 0.8100 1.5750 0.9375 ;
        RECT 1.4775 0.2625 1.5525 0.5700 ;
        RECT 1.3275 0.6450 1.5525 0.7200 ;
        RECT 1.3425 0.2625 1.4775 0.3375 ;
        RECT 0.8625 0.8625 1.4775 0.9375 ;
        RECT 1.2525 0.4125 1.3275 0.7200 ;
        RECT 1.2225 0.4125 1.2525 0.4875 ;
        RECT 1.1475 0.2625 1.2225 0.4875 ;
        RECT 1.0125 0.6375 1.1775 0.7875 ;
        RECT 0.2475 0.2625 1.1475 0.3375 ;
        RECT 0.9375 0.4125 1.0125 0.7875 ;
        RECT 0.4425 0.4125 0.9375 0.4875 ;
        RECT 0.7875 0.5625 0.8625 0.9375 ;
        RECT 0.6525 0.5625 0.7875 0.6375 ;
    END
END LHQ_1010


MACRO LNQ_0011
    CLASS CORE ;
    FOREIGN LNQ_0011 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.3100 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 2.1975 0.3075 2.2725 0.7425 ;
        RECT 2.0325 0.3075 2.1975 0.3825 ;
        RECT 2.0325 0.6675 2.1975 0.7425 ;
        RECT 1.9575 0.2100 2.0325 0.3825 ;
        RECT 1.9575 0.6675 2.0325 0.8475 ;
        END
    END Q
    PIN EN
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.2025 0.7125 0.6675 0.7875 ;
        VIA 0.3150 0.7500 VIA12_square ;
        END
    END EN
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.6275 0.1125 1.7400 0.4125 ;
        RECT 1.1625 0.1125 1.6275 0.1875 ;
        VIA 1.6875 0.3375 VIA12_square ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 2.2650 -0.0750 2.3100 0.0750 ;
        RECT 2.1450 -0.0750 2.2650 0.2325 ;
        RECT 1.8450 -0.0750 2.1450 0.0750 ;
        RECT 1.7250 -0.0750 1.8450 0.1800 ;
        RECT 1.0050 -0.0750 1.7250 0.0750 ;
        RECT 0.8850 -0.0750 1.0050 0.1800 ;
        RECT 0.3750 -0.0750 0.8850 0.0750 ;
        RECT 0.2550 -0.0750 0.3750 0.1875 ;
        RECT 0.0000 -0.0750 0.2550 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 2.2650 0.9750 2.3100 1.1250 ;
        RECT 2.1450 0.8175 2.2650 1.1250 ;
        RECT 1.8600 0.9750 2.1450 1.1250 ;
        RECT 1.7550 0.8400 1.8600 1.1250 ;
        RECT 1.0050 0.9750 1.7550 1.1250 ;
        RECT 0.8850 0.8700 1.0050 1.1250 ;
        RECT 0.3750 0.9750 0.8850 1.1250 ;
        RECT 0.2550 0.8625 0.3750 1.1250 ;
        RECT 0.0000 0.9750 0.2550 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 2.1750 0.1575 2.2350 0.2175 ;
        RECT 2.1750 0.8325 2.2350 0.8925 ;
        RECT 2.0625 0.4950 2.1225 0.5550 ;
        RECT 1.9650 0.2400 2.0250 0.3000 ;
        RECT 1.9650 0.7575 2.0250 0.8175 ;
        RECT 1.8600 0.4875 1.9200 0.5475 ;
        RECT 1.7550 0.1200 1.8150 0.1800 ;
        RECT 1.7550 0.8700 1.8150 0.9300 ;
        RECT 1.6425 0.4425 1.7025 0.5025 ;
        RECT 1.4475 0.4200 1.5075 0.4800 ;
        RECT 1.4400 0.6600 1.5000 0.7200 ;
        RECT 1.3350 0.1575 1.3950 0.2175 ;
        RECT 1.3350 0.8325 1.3950 0.8925 ;
        RECT 1.2225 0.3300 1.2825 0.3900 ;
        RECT 1.2225 0.6600 1.2825 0.7200 ;
        RECT 1.0125 0.4875 1.0725 0.5475 ;
        RECT 0.9150 0.1200 0.9750 0.1800 ;
        RECT 0.9150 0.8700 0.9750 0.9300 ;
        RECT 0.8025 0.4950 0.8625 0.5550 ;
        RECT 0.7050 0.2325 0.7650 0.2925 ;
        RECT 0.7050 0.7500 0.7650 0.8100 ;
        RECT 0.4950 0.1800 0.5550 0.2400 ;
        RECT 0.4950 0.8100 0.5550 0.8700 ;
        RECT 0.3825 0.3975 0.4425 0.4575 ;
        RECT 0.2850 0.1275 0.3450 0.1875 ;
        RECT 0.2850 0.8700 0.3450 0.9300 ;
        RECT 0.1875 0.5925 0.2475 0.6525 ;
        RECT 0.0750 0.1725 0.1350 0.2325 ;
        RECT 0.0750 0.8100 0.1350 0.8700 ;
        LAYER M1 ;
        RECT 1.8825 0.4650 2.1225 0.5850 ;
        RECT 1.8075 0.4650 1.8825 0.6825 ;
        RECT 1.7325 0.2550 1.8600 0.3675 ;
        RECT 1.6275 0.2550 1.7325 0.5400 ;
        RECT 1.4625 0.6300 1.6800 0.7200 ;
        RECT 1.5300 0.7950 1.6800 0.9000 ;
        RECT 1.3875 0.1500 1.5525 0.3450 ;
        RECT 1.4175 0.4200 1.5375 0.5550 ;
        RECT 1.2900 0.8250 1.5300 0.9000 ;
        RECT 1.3575 0.6300 1.4625 0.7500 ;
        RECT 1.2825 0.4800 1.4175 0.5550 ;
        RECT 1.2975 0.1500 1.3875 0.2250 ;
        RECT 1.1925 0.3000 1.3125 0.4050 ;
        RECT 1.2075 0.4800 1.2825 0.7500 ;
        RECT 1.1625 0.6300 1.2075 0.7500 ;
        RECT 1.0875 0.1500 1.1925 0.4050 ;
        RECT 1.0875 0.6300 1.1625 0.8325 ;
        RECT 1.0125 0.4800 1.1025 0.5550 ;
        RECT 0.9375 0.2625 1.0125 0.7950 ;
        RECT 0.7950 0.2625 0.9375 0.3375 ;
        RECT 0.7725 0.7200 0.9375 0.7950 ;
        RECT 0.6675 0.4125 0.8625 0.6450 ;
        RECT 0.7050 0.1950 0.7950 0.3375 ;
        RECT 0.6975 0.7200 0.7725 0.8700 ;
        RECT 0.5175 0.1500 0.5925 0.9000 ;
        RECT 0.4875 0.1500 0.5175 0.2700 ;
        RECT 0.4875 0.7800 0.5175 0.9000 ;
        RECT 0.3375 0.3675 0.4425 0.4875 ;
        RECT 0.2325 0.5625 0.3975 0.7875 ;
        RECT 0.1575 0.4125 0.3375 0.4875 ;
        RECT 0.1875 0.5625 0.2325 0.6825 ;
        RECT 0.1125 0.1500 0.1575 0.4875 ;
        RECT 0.1125 0.7800 0.1425 0.9000 ;
        RECT 0.0375 0.1500 0.1125 0.9000 ;
        LAYER VIA1 ;
        RECT 1.8075 0.5625 1.8825 0.6375 ;
        RECT 1.5675 0.8100 1.6425 0.8850 ;
        RECT 1.4325 0.2625 1.5075 0.3375 ;
        RECT 1.4025 0.6450 1.4775 0.7200 ;
        RECT 1.1025 0.2625 1.1775 0.3375 ;
        RECT 1.0875 0.6750 1.1625 0.7500 ;
        RECT 0.7275 0.5625 0.8025 0.6375 ;
        RECT 0.5175 0.2625 0.5925 0.3375 ;
        RECT 0.3225 0.4125 0.3975 0.4875 ;
        LAYER M2 ;
        RECT 1.7475 0.5625 1.9650 0.6375 ;
        RECT 1.6725 0.4950 1.7475 0.8850 ;
        RECT 1.5525 0.4950 1.6725 0.5700 ;
        RECT 1.5750 0.8100 1.6725 0.8850 ;
        RECT 1.4775 0.8100 1.5750 0.9375 ;
        RECT 1.4775 0.2625 1.5525 0.5700 ;
        RECT 1.3275 0.6450 1.5525 0.7200 ;
        RECT 1.3425 0.2625 1.4775 0.3375 ;
        RECT 0.8625 0.8625 1.4775 0.9375 ;
        RECT 1.2525 0.4125 1.3275 0.7200 ;
        RECT 1.2225 0.4125 1.2525 0.4875 ;
        RECT 1.1475 0.2625 1.2225 0.4875 ;
        RECT 1.0125 0.6375 1.1775 0.7875 ;
        RECT 0.4725 0.2625 1.1475 0.3375 ;
        RECT 0.9375 0.4125 1.0125 0.7875 ;
        RECT 0.2475 0.4125 0.9375 0.4875 ;
        RECT 0.7875 0.5625 0.8625 0.9375 ;
        RECT 0.6525 0.5625 0.7875 0.6375 ;
    END
END LNQ_0011


MACRO LNQ_0111
    CLASS CORE ;
    FOREIGN LNQ_0111 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.7300 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 2.0475 0.2325 2.3625 0.7350 ;
        VIA 2.2050 0.3150 VIA12_slot ;
        VIA 2.2050 0.6525 VIA12_slot ;
        END
    END Q
    PIN EN
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.2025 0.7125 0.6675 0.7875 ;
        VIA 0.3150 0.7500 VIA12_square ;
        END
    END EN
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.6275 0.1125 1.7400 0.4125 ;
        RECT 1.1625 0.1125 1.6275 0.1875 ;
        VIA 1.6875 0.3375 VIA12_square ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 2.6625 -0.0750 2.7300 0.0750 ;
        RECT 2.5875 -0.0750 2.6625 0.2475 ;
        RECT 2.2650 -0.0750 2.5875 0.0750 ;
        RECT 2.1450 -0.0750 2.2650 0.1875 ;
        RECT 1.8450 -0.0750 2.1450 0.0750 ;
        RECT 1.7250 -0.0750 1.8450 0.1800 ;
        RECT 1.0050 -0.0750 1.7250 0.0750 ;
        RECT 0.8850 -0.0750 1.0050 0.1800 ;
        RECT 0.3750 -0.0750 0.8850 0.0750 ;
        RECT 0.2550 -0.0750 0.3750 0.1875 ;
        RECT 0.0000 -0.0750 0.2550 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 2.6850 0.9750 2.7300 1.1250 ;
        RECT 2.5650 0.6450 2.6850 1.1250 ;
        RECT 2.2650 0.9750 2.5650 1.1250 ;
        RECT 2.1450 0.8175 2.2650 1.1250 ;
        RECT 1.8600 0.9750 2.1450 1.1250 ;
        RECT 1.7550 0.8400 1.8600 1.1250 ;
        RECT 1.0050 0.9750 1.7550 1.1250 ;
        RECT 0.8850 0.8700 1.0050 1.1250 ;
        RECT 0.3750 0.9750 0.8850 1.1250 ;
        RECT 0.2550 0.8625 0.3750 1.1250 ;
        RECT 0.0000 0.9750 0.2550 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 2.5950 0.1575 2.6550 0.2175 ;
        RECT 2.5950 0.6675 2.6550 0.7275 ;
        RECT 2.5950 0.8325 2.6550 0.8925 ;
        RECT 2.4900 0.4725 2.5500 0.5325 ;
        RECT 2.3850 0.2850 2.4450 0.3450 ;
        RECT 2.3850 0.6525 2.4450 0.7125 ;
        RECT 2.2800 0.4725 2.3400 0.5325 ;
        RECT 2.1750 0.1275 2.2350 0.1875 ;
        RECT 2.1750 0.8325 2.2350 0.8925 ;
        RECT 2.0700 0.4725 2.1300 0.5325 ;
        RECT 1.9650 0.2700 2.0250 0.3300 ;
        RECT 1.9650 0.6525 2.0250 0.7125 ;
        RECT 1.8600 0.4725 1.9200 0.5325 ;
        RECT 1.7550 0.1200 1.8150 0.1800 ;
        RECT 1.7550 0.8700 1.8150 0.9300 ;
        RECT 1.6425 0.4425 1.7025 0.5025 ;
        RECT 1.4475 0.4200 1.5075 0.4800 ;
        RECT 1.4400 0.6600 1.5000 0.7200 ;
        RECT 1.3350 0.1575 1.3950 0.2175 ;
        RECT 1.3350 0.8325 1.3950 0.8925 ;
        RECT 1.2225 0.3300 1.2825 0.3900 ;
        RECT 1.2225 0.6600 1.2825 0.7200 ;
        RECT 1.0125 0.4875 1.0725 0.5475 ;
        RECT 0.9150 0.1200 0.9750 0.1800 ;
        RECT 0.9150 0.8700 0.9750 0.9300 ;
        RECT 0.8025 0.4950 0.8625 0.5550 ;
        RECT 0.7050 0.2325 0.7650 0.2925 ;
        RECT 0.7050 0.7500 0.7650 0.8100 ;
        RECT 0.4950 0.1800 0.5550 0.2400 ;
        RECT 0.4950 0.8100 0.5550 0.8700 ;
        RECT 0.3825 0.3975 0.4425 0.4575 ;
        RECT 0.2850 0.1275 0.3450 0.1875 ;
        RECT 0.2850 0.8700 0.3450 0.9300 ;
        RECT 0.1875 0.5925 0.2475 0.6525 ;
        RECT 0.0750 0.1725 0.1350 0.2325 ;
        RECT 0.0750 0.8100 0.1350 0.8700 ;
        LAYER M1 ;
        RECT 1.8825 0.4650 2.5800 0.5400 ;
        RECT 2.0475 0.2625 2.4750 0.3600 ;
        RECT 1.9650 0.6150 2.4675 0.7425 ;
        RECT 1.9650 0.2400 2.0475 0.3600 ;
        RECT 1.8075 0.4650 1.8825 0.6825 ;
        RECT 1.7325 0.2550 1.8600 0.3675 ;
        RECT 1.6275 0.2550 1.7325 0.5400 ;
        RECT 1.4625 0.6300 1.6800 0.7200 ;
        RECT 1.5300 0.7950 1.6800 0.9000 ;
        RECT 1.3875 0.1500 1.5525 0.3450 ;
        RECT 1.4175 0.4200 1.5375 0.5550 ;
        RECT 1.2900 0.8250 1.5300 0.9000 ;
        RECT 1.3575 0.6300 1.4625 0.7500 ;
        RECT 1.2825 0.4800 1.4175 0.5550 ;
        RECT 1.2975 0.1500 1.3875 0.2250 ;
        RECT 1.1925 0.3000 1.3125 0.4050 ;
        RECT 1.2075 0.4800 1.2825 0.7500 ;
        RECT 1.1625 0.6300 1.2075 0.7500 ;
        RECT 1.0875 0.1500 1.1925 0.4050 ;
        RECT 1.0875 0.6300 1.1625 0.8325 ;
        RECT 1.0125 0.4800 1.1025 0.5550 ;
        RECT 0.9375 0.2625 1.0125 0.7950 ;
        RECT 0.7950 0.2625 0.9375 0.3375 ;
        RECT 0.7725 0.7200 0.9375 0.7950 ;
        RECT 0.6675 0.4125 0.8625 0.6450 ;
        RECT 0.7050 0.1950 0.7950 0.3375 ;
        RECT 0.6975 0.7200 0.7725 0.8700 ;
        RECT 0.5175 0.1500 0.5925 0.9000 ;
        RECT 0.4875 0.1500 0.5175 0.2700 ;
        RECT 0.4875 0.7800 0.5175 0.9000 ;
        RECT 0.3375 0.3675 0.4425 0.4875 ;
        RECT 0.2325 0.5625 0.3975 0.7875 ;
        RECT 0.1575 0.4125 0.3375 0.4875 ;
        RECT 0.1875 0.5625 0.2325 0.6825 ;
        RECT 0.1125 0.1500 0.1575 0.4875 ;
        RECT 0.1125 0.7800 0.1425 0.9000 ;
        RECT 0.0375 0.1500 0.1125 0.9000 ;
        LAYER VIA1 ;
        RECT 1.8075 0.5625 1.8825 0.6375 ;
        RECT 1.5675 0.8100 1.6425 0.8850 ;
        RECT 1.4325 0.2625 1.5075 0.3375 ;
        RECT 1.4025 0.6450 1.4775 0.7200 ;
        RECT 1.1025 0.2625 1.1775 0.3375 ;
        RECT 1.0875 0.6750 1.1625 0.7500 ;
        RECT 0.7275 0.5625 0.8025 0.6375 ;
        RECT 0.5175 0.2625 0.5925 0.3375 ;
        RECT 0.3225 0.4125 0.3975 0.4875 ;
        LAYER M2 ;
        RECT 1.8075 0.4950 1.8825 0.8850 ;
        RECT 1.5525 0.4950 1.8075 0.5700 ;
        RECT 1.5750 0.8100 1.8075 0.8850 ;
        RECT 1.4775 0.8100 1.5750 0.9375 ;
        RECT 1.4775 0.2625 1.5525 0.5700 ;
        RECT 1.3275 0.6450 1.5525 0.7200 ;
        RECT 1.3425 0.2625 1.4775 0.3375 ;
        RECT 0.8625 0.8625 1.4775 0.9375 ;
        RECT 1.2525 0.4125 1.3275 0.7200 ;
        RECT 1.2225 0.4125 1.2525 0.4875 ;
        RECT 1.1475 0.2625 1.2225 0.4875 ;
        RECT 1.0125 0.6375 1.1775 0.7875 ;
        RECT 0.4725 0.2625 1.1475 0.3375 ;
        RECT 0.9375 0.4125 1.0125 0.7875 ;
        RECT 0.2475 0.4125 0.9375 0.4875 ;
        RECT 0.7875 0.5625 0.8625 0.9375 ;
        RECT 0.6525 0.5625 0.7875 0.6375 ;
    END
END LNQ_0111


MACRO LNQ_1010
    CLASS CORE ;
    FOREIGN LNQ_1010 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.1000 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 1.9875 0.2175 2.0625 0.8325 ;
        RECT 1.9575 0.2175 1.9875 0.3825 ;
        RECT 1.9650 0.6675 1.9875 0.8325 ;
        END
    END Q
    PIN EN
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.2025 0.7125 0.6675 0.7875 ;
        VIA 0.3150 0.7500 VIA12_square ;
        END
    END EN
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.6275 0.1125 1.7400 0.4125 ;
        RECT 1.1625 0.1125 1.6275 0.1875 ;
        VIA 1.6875 0.3375 VIA12_square ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.8450 -0.0750 2.1000 0.0750 ;
        RECT 1.7250 -0.0750 1.8450 0.1800 ;
        RECT 1.0050 -0.0750 1.7250 0.0750 ;
        RECT 0.8850 -0.0750 1.0050 0.1800 ;
        RECT 0.3750 -0.0750 0.8850 0.0750 ;
        RECT 0.2550 -0.0750 0.3750 0.1875 ;
        RECT 0.0000 -0.0750 0.2550 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.8600 0.9750 2.1000 1.1250 ;
        RECT 1.7550 0.8400 1.8600 1.1250 ;
        RECT 1.0050 0.9750 1.7550 1.1250 ;
        RECT 0.8850 0.8700 1.0050 1.1250 ;
        RECT 0.3750 0.9750 0.8850 1.1250 ;
        RECT 0.2550 0.8625 0.3750 1.1250 ;
        RECT 0.0000 0.9750 0.2550 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.9650 0.2700 2.0250 0.3300 ;
        RECT 1.9650 0.7200 2.0250 0.7800 ;
        RECT 1.8525 0.4725 1.9125 0.5325 ;
        RECT 1.7550 0.1200 1.8150 0.1800 ;
        RECT 1.7550 0.8700 1.8150 0.9300 ;
        RECT 1.6425 0.4425 1.7025 0.5025 ;
        RECT 1.4475 0.4200 1.5075 0.4800 ;
        RECT 1.4400 0.6600 1.5000 0.7200 ;
        RECT 1.3350 0.1575 1.3950 0.2175 ;
        RECT 1.3350 0.8325 1.3950 0.8925 ;
        RECT 1.2225 0.3300 1.2825 0.3900 ;
        RECT 1.2225 0.6600 1.2825 0.7200 ;
        RECT 1.0125 0.4875 1.0725 0.5475 ;
        RECT 0.9150 0.1200 0.9750 0.1800 ;
        RECT 0.9150 0.8700 0.9750 0.9300 ;
        RECT 0.8025 0.4950 0.8625 0.5550 ;
        RECT 0.7050 0.2325 0.7650 0.2925 ;
        RECT 0.7050 0.7500 0.7650 0.8100 ;
        RECT 0.4950 0.1800 0.5550 0.2400 ;
        RECT 0.4950 0.8100 0.5550 0.8700 ;
        RECT 0.3825 0.3975 0.4425 0.4575 ;
        RECT 0.2850 0.1275 0.3450 0.1875 ;
        RECT 0.2850 0.8700 0.3450 0.9300 ;
        RECT 0.1875 0.5925 0.2475 0.6525 ;
        RECT 0.0750 0.1725 0.1350 0.2325 ;
        RECT 0.0750 0.8100 0.1350 0.8700 ;
        LAYER M1 ;
        RECT 1.8900 0.4425 1.9125 0.6075 ;
        RECT 1.8075 0.4425 1.8900 0.7650 ;
        RECT 1.7325 0.2550 1.8600 0.3675 ;
        RECT 1.7850 0.6000 1.8075 0.7650 ;
        RECT 1.6275 0.2550 1.7325 0.5400 ;
        RECT 1.4625 0.6300 1.6800 0.7200 ;
        RECT 1.5300 0.7950 1.6800 0.9000 ;
        RECT 1.3875 0.1500 1.5525 0.3450 ;
        RECT 1.4175 0.4200 1.5375 0.5550 ;
        RECT 1.2900 0.8250 1.5300 0.9000 ;
        RECT 1.3575 0.6300 1.4625 0.7500 ;
        RECT 1.2825 0.4800 1.4175 0.5550 ;
        RECT 1.2975 0.1500 1.3875 0.2250 ;
        RECT 1.1925 0.3000 1.3125 0.4050 ;
        RECT 1.2075 0.4800 1.2825 0.7500 ;
        RECT 1.1625 0.6300 1.2075 0.7500 ;
        RECT 1.0875 0.1500 1.1925 0.4050 ;
        RECT 1.0875 0.6300 1.1625 0.8325 ;
        RECT 1.0125 0.4800 1.1025 0.5550 ;
        RECT 0.9375 0.2625 1.0125 0.7950 ;
        RECT 0.7950 0.2625 0.9375 0.3375 ;
        RECT 0.7725 0.7200 0.9375 0.7950 ;
        RECT 0.6675 0.4125 0.8625 0.6450 ;
        RECT 0.7050 0.1950 0.7950 0.3375 ;
        RECT 0.6975 0.7200 0.7725 0.8700 ;
        RECT 0.5175 0.1500 0.5925 0.9000 ;
        RECT 0.4875 0.1500 0.5175 0.2700 ;
        RECT 0.4875 0.7800 0.5175 0.9000 ;
        RECT 0.3375 0.3675 0.4425 0.4875 ;
        RECT 0.2325 0.5625 0.3975 0.7875 ;
        RECT 0.1575 0.4125 0.3375 0.4875 ;
        RECT 0.1875 0.5625 0.2325 0.6825 ;
        RECT 0.1125 0.1500 0.1575 0.4875 ;
        RECT 0.1125 0.7800 0.1425 0.9000 ;
        RECT 0.0375 0.1500 0.1125 0.9000 ;
        LAYER VIA1 ;
        RECT 1.8150 0.5625 1.8900 0.6375 ;
        RECT 1.5675 0.8100 1.6425 0.8850 ;
        RECT 1.4325 0.2625 1.5075 0.3375 ;
        RECT 1.4025 0.6450 1.4775 0.7200 ;
        RECT 1.1025 0.2625 1.1775 0.3375 ;
        RECT 1.0875 0.6750 1.1625 0.7500 ;
        RECT 0.7275 0.5625 0.8025 0.6375 ;
        RECT 0.5175 0.2625 0.5925 0.3375 ;
        RECT 0.3225 0.4125 0.3975 0.4875 ;
        LAYER M2 ;
        RECT 1.7475 0.5625 1.9650 0.6375 ;
        RECT 1.6725 0.4950 1.7475 0.8850 ;
        RECT 1.5525 0.4950 1.6725 0.5700 ;
        RECT 1.5750 0.8100 1.6725 0.8850 ;
        RECT 1.4775 0.8100 1.5750 0.9375 ;
        RECT 1.4775 0.2625 1.5525 0.5700 ;
        RECT 1.3275 0.6450 1.5525 0.7200 ;
        RECT 1.3425 0.2625 1.4775 0.3375 ;
        RECT 0.8625 0.8625 1.4775 0.9375 ;
        RECT 1.2525 0.4125 1.3275 0.7200 ;
        RECT 1.2225 0.4125 1.2525 0.4875 ;
        RECT 1.1475 0.2625 1.2225 0.4875 ;
        RECT 1.0125 0.6375 1.1775 0.7875 ;
        RECT 0.4725 0.2625 1.1475 0.3375 ;
        RECT 0.9375 0.4125 1.0125 0.7875 ;
        RECT 0.2475 0.4125 0.9375 0.4875 ;
        RECT 0.7875 0.5625 0.8625 0.9375 ;
        RECT 0.6525 0.5625 0.7875 0.6375 ;
    END
END LNQ_1010


MACRO MAOI222_0011
    CLASS CORE ;
    FOREIGN MAOI222_0011 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.1000 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 1.9875 0.2925 2.0625 0.7125 ;
        RECT 1.8225 0.2925 1.9875 0.3675 ;
        RECT 1.8225 0.6375 1.9875 0.7125 ;
        RECT 1.7475 0.1950 1.8225 0.3675 ;
        RECT 1.7475 0.6375 1.8225 0.8325 ;
        END
    END ZN
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.2475 0.4125 0.7125 0.4875 ;
        VIA 0.6300 0.4500 VIA12_square ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.3525 0.5625 0.8175 0.6375 ;
        VIA 0.4350 0.6000 VIA12_square ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.0125 0.4650 1.1775 0.5400 ;
        RECT 0.9375 0.4650 1.0125 0.7875 ;
        RECT 0.1725 0.7125 0.9375 0.7875 ;
        VIA 1.0950 0.5025 VIA12_square ;
        VIA 0.2550 0.7500 VIA12_square ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 2.0550 -0.0750 2.1000 0.0750 ;
        RECT 1.9350 -0.0750 2.0550 0.2175 ;
        RECT 1.6350 -0.0750 1.9350 0.0750 ;
        RECT 1.5150 -0.0750 1.6350 0.1875 ;
        RECT 0.5850 -0.0750 1.5150 0.0750 ;
        RECT 0.4650 -0.0750 0.5850 0.1875 ;
        RECT 0.0000 -0.0750 0.4650 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 2.0475 0.9750 2.1000 1.1250 ;
        RECT 1.9425 0.8025 2.0475 1.1250 ;
        RECT 1.6350 0.9750 1.9425 1.1250 ;
        RECT 1.5150 0.8475 1.6350 1.1250 ;
        RECT 0.5625 0.9750 1.5150 1.1250 ;
        RECT 0.4575 0.8400 0.5625 1.1250 ;
        RECT 0.0000 0.9750 0.4575 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.9650 0.1575 2.0250 0.2175 ;
        RECT 1.9650 0.8325 2.0250 0.8925 ;
        RECT 1.8525 0.4725 1.9125 0.5325 ;
        RECT 1.7550 0.2250 1.8150 0.2850 ;
        RECT 1.7550 0.7200 1.8150 0.7800 ;
        RECT 1.6500 0.4725 1.7100 0.5325 ;
        RECT 1.5450 0.1275 1.6050 0.1875 ;
        RECT 1.5450 0.8550 1.6050 0.9150 ;
        RECT 1.4400 0.4650 1.5000 0.5250 ;
        RECT 1.3350 0.2250 1.3950 0.2850 ;
        RECT 1.3350 0.7575 1.3950 0.8175 ;
        RECT 1.1250 0.1575 1.1850 0.2175 ;
        RECT 1.1250 0.8325 1.1850 0.8925 ;
        RECT 1.0200 0.4875 1.0800 0.5475 ;
        RECT 0.9150 0.3000 0.9750 0.3600 ;
        RECT 0.9150 0.6675 0.9750 0.7275 ;
        RECT 0.8025 0.4950 0.8625 0.5550 ;
        RECT 0.7050 0.1575 0.7650 0.2175 ;
        RECT 0.7050 0.8325 0.7650 0.8925 ;
        RECT 0.6000 0.4800 0.6600 0.5400 ;
        RECT 0.4950 0.1200 0.5550 0.1800 ;
        RECT 0.4950 0.8700 0.5550 0.9300 ;
        RECT 0.3900 0.4800 0.4500 0.5400 ;
        RECT 0.1875 0.4800 0.2475 0.5400 ;
        RECT 0.0750 0.3000 0.1350 0.3600 ;
        RECT 0.0750 0.6750 0.1350 0.7350 ;
        LAYER M1 ;
        RECT 1.6575 0.4425 1.9125 0.5625 ;
        RECT 1.5825 0.2625 1.6575 0.7725 ;
        RECT 1.4025 0.2625 1.5825 0.3375 ;
        RECT 1.4025 0.6975 1.5825 0.7725 ;
        RECT 1.3500 0.4125 1.5000 0.6225 ;
        RECT 1.3275 0.1950 1.4025 0.3375 ;
        RECT 1.3275 0.6975 1.4025 0.8700 ;
        RECT 1.1175 0.4650 1.2750 0.5850 ;
        RECT 0.7650 0.1500 1.2225 0.2250 ;
        RECT 0.8325 0.3000 1.2225 0.3900 ;
        RECT 1.0575 0.6600 1.2225 0.7500 ;
        RECT 0.6750 0.8250 1.2150 0.9000 ;
        RECT 0.9975 0.4650 1.1175 0.5700 ;
        RECT 0.8925 0.6450 1.0575 0.7500 ;
        RECT 0.8175 0.4950 0.8925 0.5700 ;
        RECT 0.7425 0.4950 0.8175 0.7500 ;
        RECT 0.6600 0.1500 0.7650 0.2550 ;
        RECT 0.4725 0.6750 0.7425 0.7500 ;
        RECT 0.6675 0.3300 0.7200 0.4200 ;
        RECT 0.5925 0.3300 0.6675 0.6000 ;
        RECT 0.5475 0.4425 0.5925 0.6000 ;
        RECT 0.3525 0.2625 0.5175 0.3675 ;
        RECT 0.3975 0.4500 0.4725 0.7500 ;
        RECT 0.3675 0.4500 0.3975 0.5700 ;
        RECT 0.1125 0.2925 0.3525 0.3675 ;
        RECT 0.2175 0.4500 0.2925 0.8550 ;
        RECT 0.1875 0.4500 0.2175 0.5700 ;
        RECT 0.1125 0.6450 0.1350 0.7650 ;
        RECT 0.0375 0.2925 0.1125 0.7650 ;
        LAYER VIA1 ;
        RECT 1.3725 0.4650 1.4475 0.5400 ;
        RECT 1.1025 0.6750 1.1775 0.7500 ;
        RECT 0.8775 0.3000 0.9525 0.3750 ;
        RECT 0.3975 0.2625 0.4725 0.3375 ;
        LAYER M2 ;
        RECT 1.3725 0.2625 1.4475 0.7875 ;
        RECT 0.9975 0.2625 1.3725 0.3375 ;
        RECT 1.1925 0.7125 1.3725 0.7875 ;
        RECT 1.0875 0.6300 1.1925 0.7875 ;
        RECT 0.8325 0.2625 0.9975 0.3750 ;
        RECT 0.3525 0.2625 0.8325 0.3375 ;
    END
END MAOI222_0011


MACRO MAOI222_0111
    CLASS CORE ;
    FOREIGN MAOI222_0111 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.5200 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 1.8375 0.2625 2.1525 0.7500 ;
        VIA 1.9950 0.3450 VIA12_slot ;
        VIA 1.9950 0.6675 VIA12_slot ;
        END
    END ZN
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.2475 0.4125 0.7125 0.4875 ;
        VIA 0.6300 0.4500 VIA12_square ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.3525 0.5625 0.8175 0.6375 ;
        VIA 0.4350 0.6000 VIA12_square ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.0125 0.4650 1.1775 0.5400 ;
        RECT 0.9375 0.4650 1.0125 0.7875 ;
        RECT 0.1725 0.7125 0.9375 0.7875 ;
        VIA 1.0950 0.5025 VIA12_square ;
        VIA 0.2550 0.7500 VIA12_square ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 2.4525 -0.0750 2.5200 0.0750 ;
        RECT 2.3775 -0.0750 2.4525 0.3150 ;
        RECT 2.0550 -0.0750 2.3775 0.0750 ;
        RECT 1.9350 -0.0750 2.0550 0.1950 ;
        RECT 1.6350 -0.0750 1.9350 0.0750 ;
        RECT 1.5150 -0.0750 1.6350 0.1875 ;
        RECT 0.5850 -0.0750 1.5150 0.0750 ;
        RECT 0.4650 -0.0750 0.5850 0.1875 ;
        RECT 0.0000 -0.0750 0.4650 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 2.4525 0.9750 2.5200 1.1250 ;
        RECT 2.3775 0.6375 2.4525 1.1250 ;
        RECT 2.0325 0.9750 2.3775 1.1250 ;
        RECT 1.9575 0.8175 2.0325 1.1250 ;
        RECT 1.6350 0.9750 1.9575 1.1250 ;
        RECT 1.5150 0.8475 1.6350 1.1250 ;
        RECT 0.5625 0.9750 1.5150 1.1250 ;
        RECT 0.4575 0.8400 0.5625 1.1250 ;
        RECT 0.0000 0.9750 0.4575 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 2.3850 0.2250 2.4450 0.2850 ;
        RECT 2.3850 0.6675 2.4450 0.7275 ;
        RECT 2.3850 0.8325 2.4450 0.8925 ;
        RECT 2.2800 0.4650 2.3400 0.5250 ;
        RECT 2.1750 0.2250 2.2350 0.2850 ;
        RECT 2.1750 0.7200 2.2350 0.7800 ;
        RECT 2.0700 0.4650 2.1300 0.5250 ;
        RECT 1.9650 0.1275 2.0250 0.1875 ;
        RECT 1.9650 0.8475 2.0250 0.9075 ;
        RECT 1.8600 0.4650 1.9200 0.5250 ;
        RECT 1.7550 0.2250 1.8150 0.2850 ;
        RECT 1.7550 0.7200 1.8150 0.7800 ;
        RECT 1.6500 0.4725 1.7100 0.5325 ;
        RECT 1.5450 0.1275 1.6050 0.1875 ;
        RECT 1.5450 0.8550 1.6050 0.9150 ;
        RECT 1.4400 0.4650 1.5000 0.5250 ;
        RECT 1.3350 0.2250 1.3950 0.2850 ;
        RECT 1.3350 0.7575 1.3950 0.8175 ;
        RECT 1.1250 0.1575 1.1850 0.2175 ;
        RECT 1.1250 0.8325 1.1850 0.8925 ;
        RECT 1.0200 0.4875 1.0800 0.5475 ;
        RECT 0.9150 0.3000 0.9750 0.3600 ;
        RECT 0.9150 0.6675 0.9750 0.7275 ;
        RECT 0.8025 0.4950 0.8625 0.5550 ;
        RECT 0.7050 0.1575 0.7650 0.2175 ;
        RECT 0.7050 0.8325 0.7650 0.8925 ;
        RECT 0.6000 0.4800 0.6600 0.5400 ;
        RECT 0.4950 0.1200 0.5550 0.1800 ;
        RECT 0.4950 0.8700 0.5550 0.9300 ;
        RECT 0.3900 0.4800 0.4500 0.5400 ;
        RECT 0.1875 0.4800 0.2475 0.5400 ;
        RECT 0.0750 0.3000 0.1350 0.3600 ;
        RECT 0.0750 0.6750 0.1350 0.7350 ;
        LAYER M1 ;
        RECT 1.6575 0.4575 2.3700 0.5325 ;
        RECT 2.1525 0.1950 2.2575 0.3825 ;
        RECT 2.1675 0.6225 2.2425 0.8325 ;
        RECT 1.8225 0.6225 2.1675 0.7125 ;
        RECT 1.8375 0.2925 2.1525 0.3825 ;
        RECT 1.7325 0.1950 1.8375 0.3825 ;
        RECT 1.7475 0.6225 1.8225 0.8325 ;
        RECT 1.5825 0.2625 1.6575 0.7725 ;
        RECT 1.4025 0.2625 1.5825 0.3375 ;
        RECT 1.4025 0.6975 1.5825 0.7725 ;
        RECT 1.3500 0.4125 1.5000 0.6225 ;
        RECT 1.3275 0.1950 1.4025 0.3375 ;
        RECT 1.3275 0.6975 1.4025 0.8700 ;
        RECT 1.1175 0.4650 1.2750 0.5850 ;
        RECT 0.7650 0.1500 1.2225 0.2250 ;
        RECT 0.8325 0.3000 1.2225 0.3900 ;
        RECT 1.0575 0.6600 1.2225 0.7500 ;
        RECT 0.6750 0.8250 1.2150 0.9000 ;
        RECT 0.9975 0.4650 1.1175 0.5700 ;
        RECT 0.8925 0.6450 1.0575 0.7500 ;
        RECT 0.8175 0.4950 0.8925 0.5700 ;
        RECT 0.7425 0.4950 0.8175 0.7500 ;
        RECT 0.6600 0.1500 0.7650 0.2550 ;
        RECT 0.4725 0.6750 0.7425 0.7500 ;
        RECT 0.6675 0.3300 0.7200 0.4200 ;
        RECT 0.5925 0.3300 0.6675 0.6000 ;
        RECT 0.5475 0.4425 0.5925 0.6000 ;
        RECT 0.3525 0.2625 0.5175 0.3675 ;
        RECT 0.3975 0.4500 0.4725 0.7500 ;
        RECT 0.3675 0.4500 0.3975 0.5700 ;
        RECT 0.1125 0.2925 0.3525 0.3675 ;
        RECT 0.2175 0.4500 0.2925 0.8550 ;
        RECT 0.1875 0.4500 0.2175 0.5700 ;
        RECT 0.1125 0.6450 0.1350 0.7650 ;
        RECT 0.0375 0.2925 0.1125 0.7650 ;
        LAYER VIA1 ;
        RECT 1.3725 0.4650 1.4475 0.5400 ;
        RECT 1.1025 0.6750 1.1775 0.7500 ;
        RECT 0.8775 0.3000 0.9525 0.3750 ;
        RECT 0.3975 0.2625 0.4725 0.3375 ;
        LAYER M2 ;
        RECT 1.3725 0.2625 1.4475 0.7875 ;
        RECT 0.9975 0.2625 1.3725 0.3375 ;
        RECT 1.1925 0.7125 1.3725 0.7875 ;
        RECT 1.0875 0.6300 1.1925 0.7875 ;
        RECT 0.8325 0.2625 0.9975 0.3750 ;
        RECT 0.3525 0.2625 0.8325 0.3375 ;
    END
END MAOI222_0111


MACRO MAOI222_1000
    CLASS CORE ;
    FOREIGN MAOI222_1000 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.4700 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 0.8625 0.2625 0.9675 0.4125 ;
        RECT 0.3525 0.2625 0.8625 0.3375 ;
        VIA 0.9150 0.3375 VIA12_square ;
        VIA 0.4350 0.3000 VIA12_square ;
        END
    END ZN
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.2475 0.4125 0.7125 0.4875 ;
        VIA 0.6300 0.4500 VIA12_square ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.3525 0.5625 0.8175 0.6375 ;
        VIA 0.4350 0.6000 VIA12_square ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.0425 0.4050 1.1175 0.7875 ;
        RECT 0.1875 0.7125 1.0425 0.7875 ;
        VIA 1.0800 0.5175 VIA12_square ;
        VIA 0.2700 0.7500 VIA12_square ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.5850 -0.0750 1.4700 0.0750 ;
        RECT 0.4650 -0.0750 0.5850 0.1875 ;
        RECT 0.0000 -0.0750 0.4650 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.5625 0.9750 1.4700 1.1250 ;
        RECT 0.4575 0.8400 0.5625 1.1250 ;
        RECT 0.0000 0.9750 0.4575 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.3350 0.1800 1.3950 0.2400 ;
        RECT 1.3350 0.8325 1.3950 0.8925 ;
        RECT 1.2225 0.4800 1.2825 0.5400 ;
        RECT 1.1250 0.1575 1.1850 0.2175 ;
        RECT 1.1250 0.6600 1.1850 0.7200 ;
        RECT 0.9150 0.3000 0.9750 0.3600 ;
        RECT 0.9150 0.6675 0.9750 0.7275 ;
        RECT 0.8025 0.4950 0.8625 0.5550 ;
        RECT 0.7050 0.1575 0.7650 0.2175 ;
        RECT 0.7050 0.8325 0.7650 0.8925 ;
        RECT 0.6000 0.4800 0.6600 0.5400 ;
        RECT 0.4950 0.1200 0.5550 0.1800 ;
        RECT 0.4950 0.8700 0.5550 0.9300 ;
        RECT 0.3900 0.5025 0.4500 0.5625 ;
        RECT 0.1875 0.4800 0.2475 0.5400 ;
        RECT 0.0750 0.1575 0.1350 0.2175 ;
        RECT 0.0750 0.8175 0.1350 0.8775 ;
        LAYER M1 ;
        RECT 1.3575 0.1500 1.4325 0.7200 ;
        RECT 1.3200 0.7950 1.4250 0.9000 ;
        RECT 1.3200 0.1500 1.3575 0.3750 ;
        RECT 0.9975 0.6450 1.3575 0.7200 ;
        RECT 0.8325 0.3000 1.3200 0.3750 ;
        RECT 0.6750 0.8250 1.3200 0.9000 ;
        RECT 0.9975 0.4500 1.2825 0.5700 ;
        RECT 0.7650 0.1500 1.2150 0.2250 ;
        RECT 0.8925 0.6450 0.9975 0.7500 ;
        RECT 0.8175 0.4950 0.8925 0.5700 ;
        RECT 0.7425 0.4950 0.8175 0.7500 ;
        RECT 0.6600 0.1500 0.7650 0.2550 ;
        RECT 0.4725 0.6750 0.7425 0.7500 ;
        RECT 0.6675 0.3300 0.7200 0.4200 ;
        RECT 0.5925 0.3300 0.6675 0.6000 ;
        RECT 0.5475 0.4425 0.5925 0.6000 ;
        RECT 0.3525 0.2625 0.5175 0.3675 ;
        RECT 0.3975 0.4725 0.4725 0.7500 ;
        RECT 0.3825 0.4725 0.3975 0.5925 ;
        RECT 0.1650 0.2925 0.3525 0.3675 ;
        RECT 0.2325 0.4500 0.3075 0.8550 ;
        RECT 0.1875 0.4500 0.2325 0.5700 ;
        RECT 0.1125 0.1575 0.1650 0.3675 ;
        RECT 0.1125 0.7950 0.1575 0.9000 ;
        RECT 0.0375 0.1575 0.1125 0.9000 ;
    END
END MAOI222_1000


MACRO MAOI222_1010
    CLASS CORE ;
    FOREIGN MAOI222_1010 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.4700 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 0.8325 0.2625 0.9975 0.3750 ;
        RECT 0.3525 0.2625 0.8325 0.3375 ;
        VIA 0.9150 0.3375 VIA12_square ;
        VIA 0.4350 0.3000 VIA12_square ;
        END
    END ZN
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.2475 0.4125 0.7125 0.4875 ;
        VIA 0.6300 0.4500 VIA12_square ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.3525 0.5625 0.8175 0.6375 ;
        VIA 0.4350 0.6000 VIA12_square ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.0425 0.4500 1.1175 0.7875 ;
        RECT 0.1725 0.7125 1.0425 0.7875 ;
        VIA 1.0800 0.5325 VIA12_square ;
        VIA 0.2550 0.7500 VIA12_square ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.5850 -0.0750 1.4700 0.0750 ;
        RECT 0.4650 -0.0750 0.5850 0.1875 ;
        RECT 0.0000 -0.0750 0.4650 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.5625 0.9750 1.4700 1.1250 ;
        RECT 0.4575 0.8400 0.5625 1.1250 ;
        RECT 0.0000 0.9750 0.4575 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.3350 0.3000 1.3950 0.3600 ;
        RECT 1.3350 0.8325 1.3950 0.8925 ;
        RECT 1.2225 0.4800 1.2825 0.5400 ;
        RECT 1.1250 0.1575 1.1850 0.2175 ;
        RECT 1.1250 0.6600 1.1850 0.7200 ;
        RECT 0.9150 0.3000 0.9750 0.3600 ;
        RECT 0.9150 0.6675 0.9750 0.7275 ;
        RECT 0.8025 0.4950 0.8625 0.5550 ;
        RECT 0.7050 0.1575 0.7650 0.2175 ;
        RECT 0.7050 0.8325 0.7650 0.8925 ;
        RECT 0.6000 0.4800 0.6600 0.5400 ;
        RECT 0.4950 0.1200 0.5550 0.1800 ;
        RECT 0.4950 0.8700 0.5550 0.9300 ;
        RECT 0.3900 0.4800 0.4500 0.5400 ;
        RECT 0.1875 0.4800 0.2475 0.5400 ;
        RECT 0.0750 0.3000 0.1350 0.3600 ;
        RECT 0.0750 0.6750 0.1350 0.7350 ;
        LAYER M1 ;
        RECT 1.3575 0.3000 1.4325 0.7200 ;
        RECT 1.3200 0.7950 1.4250 0.9000 ;
        RECT 0.8325 0.3000 1.3575 0.3750 ;
        RECT 0.9975 0.6450 1.3575 0.7200 ;
        RECT 0.6750 0.8250 1.3200 0.9000 ;
        RECT 0.9975 0.4500 1.2825 0.5700 ;
        RECT 0.7650 0.1500 1.2225 0.2250 ;
        RECT 0.8925 0.6450 0.9975 0.7500 ;
        RECT 0.8175 0.4950 0.8925 0.5700 ;
        RECT 0.7425 0.4950 0.8175 0.7500 ;
        RECT 0.6600 0.1500 0.7650 0.2550 ;
        RECT 0.4725 0.6750 0.7425 0.7500 ;
        RECT 0.6675 0.3300 0.7200 0.4200 ;
        RECT 0.5925 0.3300 0.6675 0.6000 ;
        RECT 0.5475 0.4425 0.5925 0.6000 ;
        RECT 0.3525 0.2625 0.5175 0.3675 ;
        RECT 0.3975 0.4500 0.4725 0.7500 ;
        RECT 0.3675 0.4500 0.3975 0.5700 ;
        RECT 0.1125 0.2925 0.3525 0.3675 ;
        RECT 0.2175 0.4500 0.2925 0.8550 ;
        RECT 0.1875 0.4500 0.2175 0.5700 ;
        RECT 0.1125 0.6450 0.1350 0.7650 ;
        RECT 0.0375 0.2925 0.1125 0.7650 ;
    END
END MAOI222_1010


MACRO MAOI22_0011
    CLASS CORE ;
    FOREIGN MAOI22_0011 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.6800 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 0.9975 0.6525 1.0950 0.7575 ;
        RECT 0.9225 0.2625 0.9975 0.7575 ;
        RECT 0.5325 0.2625 0.9225 0.3375 ;
        VIA 1.0200 0.7050 VIA12_square ;
        VIA 0.9600 0.3450 VIA12_square ;
        END
    END ZN
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1425 0.4500 0.2325 0.5700 ;
        RECT 0.0675 0.3675 0.1425 0.6825 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.1875 0.7125 0.6525 0.7875 ;
        VIA 0.3450 0.7500 VIA12_square ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.1175 0.4125 1.5825 0.4875 ;
        VIA 1.2600 0.4500 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.1175 0.2625 1.5825 0.3375 ;
        VIA 1.4250 0.3000 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.2150 -0.0750 1.6800 0.0750 ;
        RECT 1.0950 -0.0750 1.2150 0.1800 ;
        RECT 0.7950 -0.0750 1.0950 0.0750 ;
        RECT 0.6900 -0.0750 0.7950 0.2250 ;
        RECT 0.0000 -0.0750 0.6900 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.6275 0.9750 1.6800 1.1250 ;
        RECT 1.5225 0.8025 1.6275 1.1250 ;
        RECT 1.2150 0.9750 1.5225 1.1250 ;
        RECT 1.0950 0.8625 1.2150 1.1250 ;
        RECT 0.7950 0.9750 1.0950 1.1250 ;
        RECT 0.6750 0.8700 0.7950 1.1250 ;
        RECT 0.1425 0.9750 0.6750 1.1250 ;
        RECT 0.0675 0.8025 0.1425 1.1250 ;
        RECT 0.0000 0.9750 0.0675 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.5450 0.2100 1.6050 0.2700 ;
        RECT 1.5450 0.8325 1.6050 0.8925 ;
        RECT 1.4325 0.4800 1.4925 0.5400 ;
        RECT 1.3350 0.6600 1.3950 0.7200 ;
        RECT 1.2300 0.4725 1.2900 0.5325 ;
        RECT 1.1250 0.1200 1.1850 0.1800 ;
        RECT 1.1250 0.8700 1.1850 0.9300 ;
        RECT 1.0125 0.4950 1.0725 0.5550 ;
        RECT 0.9150 0.2475 0.9750 0.3075 ;
        RECT 0.9150 0.6825 0.9750 0.7425 ;
        RECT 0.8100 0.4950 0.8700 0.5550 ;
        RECT 0.7050 0.1350 0.7650 0.1950 ;
        RECT 0.7050 0.8700 0.7650 0.9300 ;
        RECT 0.6000 0.4950 0.6600 0.5550 ;
        RECT 0.4950 0.1575 0.5550 0.2175 ;
        RECT 0.4950 0.7575 0.5550 0.8175 ;
        RECT 0.3825 0.4950 0.4425 0.5550 ;
        RECT 0.2850 0.3075 0.3450 0.3675 ;
        RECT 0.1725 0.4800 0.2325 0.5400 ;
        RECT 0.0750 0.1725 0.1350 0.2325 ;
        RECT 0.0750 0.8325 0.1350 0.8925 ;
        LAYER M1 ;
        RECT 1.5675 0.1800 1.6425 0.7275 ;
        RECT 1.5375 0.1800 1.5675 0.3075 ;
        RECT 1.3350 0.6525 1.5675 0.7275 ;
        RECT 1.4625 0.3900 1.4925 0.5700 ;
        RECT 1.3875 0.2175 1.4625 0.5700 ;
        RECT 1.1775 0.6525 1.3350 0.7875 ;
        RECT 1.2075 0.2550 1.3125 0.5775 ;
        RECT 0.8325 0.4950 1.1025 0.5700 ;
        RECT 1.0200 0.6525 1.1025 0.7800 ;
        RECT 1.0200 0.2475 1.0575 0.4200 ;
        RECT 0.9075 0.1500 1.0200 0.4200 ;
        RECT 0.9150 0.6525 1.0200 0.9000 ;
        RECT 0.7575 0.3000 0.8325 0.7950 ;
        RECT 0.2550 0.3000 0.7575 0.3750 ;
        RECT 0.5775 0.7200 0.7575 0.7950 ;
        RECT 0.5175 0.4500 0.6825 0.6450 ;
        RECT 0.1575 0.1500 0.5850 0.2250 ;
        RECT 0.4725 0.7200 0.5775 0.8400 ;
        RECT 0.3825 0.4500 0.4425 0.5850 ;
        RECT 0.3075 0.4500 0.3825 0.8325 ;
        RECT 0.0525 0.1500 0.1575 0.2550 ;
        LAYER VIA1 ;
        RECT 1.2150 0.6900 1.2900 0.7650 ;
        RECT 0.5625 0.5625 0.6375 0.6375 ;
        LAYER M2 ;
        RECT 1.2000 0.6525 1.3050 0.9150 ;
        RECT 0.8475 0.8400 1.2000 0.9150 ;
        RECT 0.7725 0.5625 0.8475 0.9150 ;
        RECT 0.5175 0.5625 0.7725 0.6375 ;
    END
END MAOI22_0011


MACRO MAOI22_0100
    CLASS CORE ;
    FOREIGN MAOI22_0100 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.0900 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 1.7400 0.2700 2.0550 0.7875 ;
        VIA 1.8975 0.3525 VIA12_slot ;
        VIA 1.8975 0.7050 VIA12_slot ;
        END
    END ZN
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 5.9475 0.3600 6.0225 0.6450 ;
        RECT 5.8575 0.4800 5.9475 0.6450 ;
        RECT 4.7700 0.4800 5.8575 0.5850 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 4.0950 0.5625 4.4550 0.6375 ;
        RECT 3.9900 0.4125 4.0950 0.6375 ;
        VIA 4.0425 0.5250 VIA12_square ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.2775 0.4350 1.2825 0.5625 ;
        RECT 0.1425 0.4050 0.2775 0.5625 ;
        RECT 0.0675 0.4050 0.1425 0.6825 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.4850 0.4125 1.5900 0.6000 ;
        RECT 1.0650 0.4125 1.4850 0.4875 ;
        VIA 1.5375 0.5175 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 6.0375 -0.0750 6.0900 0.0750 ;
        RECT 5.9325 -0.0750 6.0375 0.2400 ;
        RECT 5.6250 -0.0750 5.9325 0.0750 ;
        RECT 5.5050 -0.0750 5.6250 0.2175 ;
        RECT 5.2050 -0.0750 5.5050 0.0750 ;
        RECT 5.0850 -0.0750 5.2050 0.2175 ;
        RECT 4.7850 -0.0750 5.0850 0.0750 ;
        RECT 4.6650 -0.0750 4.7850 0.2175 ;
        RECT 4.3650 -0.0750 4.6650 0.0750 ;
        RECT 4.2450 -0.0750 4.3650 0.1800 ;
        RECT 3.9450 -0.0750 4.2450 0.0750 ;
        RECT 3.8250 -0.0750 3.9450 0.2175 ;
        RECT 3.3075 -0.0750 3.8250 0.0750 ;
        RECT 3.2025 -0.0750 3.3075 0.2250 ;
        RECT 2.8875 -0.0750 3.2025 0.0750 ;
        RECT 2.7825 -0.0750 2.8875 0.2250 ;
        RECT 1.2150 -0.0750 2.7825 0.0750 ;
        RECT 1.0950 -0.0750 1.2150 0.1800 ;
        RECT 0.7950 -0.0750 1.0950 0.0750 ;
        RECT 0.6750 -0.0750 0.7950 0.1800 ;
        RECT 0.3750 -0.0750 0.6750 0.0750 ;
        RECT 0.2550 -0.0750 0.3750 0.1800 ;
        RECT 0.0000 -0.0750 0.2550 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 5.8350 0.9750 6.0900 1.1250 ;
        RECT 5.7150 0.8700 5.8350 1.1250 ;
        RECT 5.4150 0.9750 5.7150 1.1250 ;
        RECT 5.2950 0.8700 5.4150 1.1250 ;
        RECT 4.9950 0.9750 5.2950 1.1250 ;
        RECT 4.8750 0.8700 4.9950 1.1250 ;
        RECT 3.3075 0.9750 4.8750 1.1250 ;
        RECT 3.2025 0.8250 3.3075 1.1250 ;
        RECT 2.8875 0.9750 3.2025 1.1250 ;
        RECT 2.7825 0.8250 2.8875 1.1250 ;
        RECT 2.4675 0.9750 2.7825 1.1250 ;
        RECT 2.3625 0.8250 2.4675 1.1250 ;
        RECT 0.0000 0.9750 2.3625 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 5.9550 0.1575 6.0150 0.2175 ;
        RECT 5.9550 0.7500 6.0150 0.8100 ;
        RECT 5.8500 0.4950 5.9100 0.5550 ;
        RECT 5.7450 0.2400 5.8050 0.3000 ;
        RECT 5.7450 0.8700 5.8050 0.9300 ;
        RECT 5.6400 0.4950 5.7000 0.5550 ;
        RECT 5.5350 0.1575 5.5950 0.2175 ;
        RECT 5.5350 0.7050 5.5950 0.7650 ;
        RECT 5.4300 0.4950 5.4900 0.5550 ;
        RECT 5.3250 0.2400 5.3850 0.3000 ;
        RECT 5.3250 0.8700 5.3850 0.9300 ;
        RECT 5.2200 0.4950 5.2800 0.5550 ;
        RECT 5.1150 0.1575 5.1750 0.2175 ;
        RECT 5.1150 0.6825 5.1750 0.7425 ;
        RECT 5.0100 0.4950 5.0700 0.5550 ;
        RECT 4.9050 0.8700 4.9650 0.9300 ;
        RECT 4.8000 0.4950 4.8600 0.5550 ;
        RECT 4.6950 0.1575 4.7550 0.2175 ;
        RECT 4.6950 0.7650 4.7550 0.8250 ;
        RECT 4.5900 0.4950 4.6500 0.5550 ;
        RECT 4.4850 0.2400 4.5450 0.3000 ;
        RECT 4.4850 0.6825 4.5450 0.7425 ;
        RECT 4.3800 0.4950 4.4400 0.5550 ;
        RECT 4.2750 0.1200 4.3350 0.1800 ;
        RECT 4.2750 0.8325 4.3350 0.8925 ;
        RECT 4.1700 0.4950 4.2300 0.5550 ;
        RECT 4.0650 0.2625 4.1250 0.3225 ;
        RECT 4.0650 0.6825 4.1250 0.7425 ;
        RECT 3.9600 0.4950 4.0200 0.5550 ;
        RECT 3.8550 0.1575 3.9150 0.2175 ;
        RECT 3.8550 0.8325 3.9150 0.8925 ;
        RECT 3.7500 0.4950 3.8100 0.5550 ;
        RECT 3.6450 0.6825 3.7050 0.7425 ;
        RECT 3.4350 0.2625 3.4950 0.3225 ;
        RECT 3.4350 0.7125 3.4950 0.7725 ;
        RECT 3.3300 0.4950 3.3900 0.5550 ;
        RECT 3.2250 0.1425 3.2850 0.2025 ;
        RECT 3.2250 0.8475 3.2850 0.9075 ;
        RECT 3.1200 0.4950 3.1800 0.5550 ;
        RECT 3.0150 0.3000 3.0750 0.3600 ;
        RECT 3.0150 0.6825 3.0750 0.7425 ;
        RECT 2.9100 0.4950 2.9700 0.5550 ;
        RECT 2.8050 0.1425 2.8650 0.2025 ;
        RECT 2.8050 0.8475 2.8650 0.9075 ;
        RECT 2.7000 0.4950 2.7600 0.5550 ;
        RECT 2.5950 0.3000 2.6550 0.3600 ;
        RECT 2.5950 0.6825 2.6550 0.7425 ;
        RECT 2.4900 0.4950 2.5500 0.5550 ;
        RECT 2.3850 0.8475 2.4450 0.9075 ;
        RECT 2.2800 0.4950 2.3400 0.5550 ;
        RECT 2.1750 0.1575 2.2350 0.2175 ;
        RECT 2.1750 0.7500 2.2350 0.8100 ;
        RECT 2.0625 0.4950 2.1225 0.5550 ;
        RECT 1.9650 0.3000 2.0250 0.3600 ;
        RECT 1.9650 0.6825 2.0250 0.7425 ;
        RECT 1.8600 0.4950 1.9200 0.5550 ;
        RECT 1.7550 0.1575 1.8150 0.2175 ;
        RECT 1.7550 0.8325 1.8150 0.8925 ;
        RECT 1.6500 0.4950 1.7100 0.5550 ;
        RECT 1.5450 0.3000 1.6050 0.3600 ;
        RECT 1.5450 0.6825 1.6050 0.7425 ;
        RECT 1.4400 0.4950 1.5000 0.5550 ;
        RECT 1.3350 0.2325 1.3950 0.2925 ;
        RECT 1.3350 0.8325 1.3950 0.8925 ;
        RECT 1.2225 0.4650 1.2825 0.5250 ;
        RECT 1.1250 0.1200 1.1850 0.1800 ;
        RECT 1.1250 0.6675 1.1850 0.7275 ;
        RECT 1.0200 0.4650 1.0800 0.5250 ;
        RECT 0.9150 0.2625 0.9750 0.3225 ;
        RECT 0.9150 0.8325 0.9750 0.8925 ;
        RECT 0.8100 0.4650 0.8700 0.5250 ;
        RECT 0.7050 0.1200 0.7650 0.1800 ;
        RECT 0.6000 0.4650 0.6600 0.5250 ;
        RECT 0.4950 0.2625 0.5550 0.3225 ;
        RECT 0.4950 0.8325 0.5550 0.8925 ;
        RECT 0.3900 0.4650 0.4500 0.5250 ;
        RECT 0.2850 0.1200 0.3450 0.1800 ;
        RECT 0.2850 0.6675 0.3450 0.7275 ;
        RECT 0.1800 0.4650 0.2400 0.5250 ;
        RECT 0.0750 0.2325 0.1350 0.2925 ;
        RECT 0.0750 0.8175 0.1350 0.8775 ;
        LAYER M1 ;
        RECT 5.9475 0.7200 6.0225 0.8400 ;
        RECT 5.6025 0.7200 5.9475 0.7950 ;
        RECT 5.7375 0.2025 5.8125 0.4050 ;
        RECT 5.3925 0.2925 5.7375 0.4050 ;
        RECT 5.5275 0.6750 5.6025 0.7950 ;
        RECT 4.7625 0.6750 5.5275 0.7500 ;
        RECT 5.3175 0.2025 5.3925 0.4050 ;
        RECT 4.5525 0.2925 5.3175 0.4050 ;
        RECT 4.6875 0.6750 4.7625 0.9000 ;
        RECT 3.8100 0.8250 4.6875 0.9000 ;
        RECT 3.7200 0.4800 4.6800 0.5850 ;
        RECT 3.6450 0.6750 4.5825 0.7500 ;
        RECT 4.4775 0.2025 4.5525 0.4050 ;
        RECT 4.1325 0.2925 4.4775 0.4050 ;
        RECT 4.0575 0.2025 4.1325 0.4050 ;
        RECT 3.6450 0.3000 4.0575 0.4050 ;
        RECT 3.5700 0.3000 3.6450 0.7500 ;
        RECT 2.2425 0.4800 3.5700 0.5850 ;
        RECT 3.4200 0.2250 3.4950 0.4050 ;
        RECT 3.4200 0.6750 3.4950 0.8100 ;
        RECT 1.5150 0.3000 3.4200 0.4050 ;
        RECT 2.2425 0.6750 3.4200 0.7500 ;
        RECT 1.4025 0.1500 2.2800 0.2250 ;
        RECT 2.1675 0.6750 2.2425 0.9000 ;
        RECT 0.1575 0.8250 2.1675 0.9000 ;
        RECT 1.3950 0.4800 2.1525 0.5850 ;
        RECT 0.2475 0.6600 2.0625 0.7500 ;
        RECT 1.3275 0.1500 1.4025 0.3300 ;
        RECT 0.1425 0.2550 1.3275 0.3300 ;
        RECT 0.0525 0.7950 0.1575 0.9000 ;
        RECT 0.0675 0.2025 0.1425 0.3300 ;
    END
END MAOI22_0100


MACRO MAOI22_0111
    CLASS CORE ;
    FOREIGN MAOI22_0111 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.1000 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 0.9975 0.2700 1.3125 0.7800 ;
        VIA 1.1550 0.3525 VIA12_slot ;
        VIA 1.1550 0.6975 VIA12_slot ;
        END
    END ZN
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1425 0.4500 0.2325 0.5700 ;
        RECT 0.0675 0.3675 0.1425 0.6825 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.4275 0.8625 0.6675 0.9375 ;
        RECT 0.3525 0.4800 0.4275 0.9375 ;
        RECT 0.1275 0.8625 0.3525 0.9375 ;
        VIA 0.3900 0.5625 VIA12_square ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.7475 0.8625 2.0250 0.9375 ;
        RECT 1.6725 0.4125 1.7475 0.9375 ;
        RECT 1.6425 0.4125 1.6725 0.5625 ;
        RECT 1.4700 0.8625 1.6725 0.9375 ;
        VIA 1.6950 0.4875 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.9575 0.3675 2.0325 0.6825 ;
        RECT 1.8600 0.4500 1.9575 0.5700 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.6350 -0.0750 2.1000 0.0750 ;
        RECT 1.5150 -0.0750 1.6350 0.1800 ;
        RECT 1.2150 -0.0750 1.5150 0.0750 ;
        RECT 1.0950 -0.0750 1.2150 0.2025 ;
        RECT 0.7950 -0.0750 1.0950 0.0750 ;
        RECT 0.6900 -0.0750 0.7950 0.2100 ;
        RECT 0.0000 -0.0750 0.6900 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 2.0325 0.9750 2.1000 1.1250 ;
        RECT 1.9575 0.8025 2.0325 1.1250 ;
        RECT 1.6350 0.9750 1.9575 1.1250 ;
        RECT 1.5150 0.8625 1.6350 1.1250 ;
        RECT 1.2150 0.9750 1.5150 1.1250 ;
        RECT 1.0950 0.8475 1.2150 1.1250 ;
        RECT 0.7950 0.9750 1.0950 1.1250 ;
        RECT 0.6750 0.8700 0.7950 1.1250 ;
        RECT 0.1425 0.9750 0.6750 1.1250 ;
        RECT 0.0675 0.8025 0.1425 1.1250 ;
        RECT 0.0000 0.9750 0.0675 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.9650 0.1725 2.0250 0.2325 ;
        RECT 1.9650 0.8325 2.0250 0.8925 ;
        RECT 1.8600 0.4800 1.9200 0.5400 ;
        RECT 1.7550 0.7275 1.8150 0.7875 ;
        RECT 1.6500 0.4800 1.7100 0.5400 ;
        RECT 1.5450 0.1200 1.6050 0.1800 ;
        RECT 1.5450 0.8700 1.6050 0.9300 ;
        RECT 1.4400 0.4950 1.5000 0.5550 ;
        RECT 1.3350 0.3075 1.3950 0.3675 ;
        RECT 1.3350 0.6825 1.3950 0.7425 ;
        RECT 1.2300 0.4950 1.2900 0.5550 ;
        RECT 1.1250 0.1350 1.1850 0.1950 ;
        RECT 1.1250 0.8550 1.1850 0.9150 ;
        RECT 1.0200 0.4950 1.0800 0.5550 ;
        RECT 0.9150 0.3075 0.9750 0.3675 ;
        RECT 0.9150 0.6825 0.9750 0.7425 ;
        RECT 0.8100 0.4950 0.8700 0.5550 ;
        RECT 0.7050 0.1200 0.7650 0.1800 ;
        RECT 0.7050 0.8700 0.7650 0.9300 ;
        RECT 0.6000 0.4950 0.6600 0.5550 ;
        RECT 0.4950 0.1575 0.5550 0.2175 ;
        RECT 0.4950 0.7575 0.5550 0.8175 ;
        RECT 0.3900 0.4950 0.4500 0.5550 ;
        RECT 0.2850 0.3075 0.3450 0.3675 ;
        RECT 0.1725 0.4800 0.2325 0.5400 ;
        RECT 0.0750 0.1725 0.1350 0.2325 ;
        RECT 0.0750 0.8325 0.1350 0.8925 ;
        LAYER M1 ;
        RECT 1.9425 0.1500 2.0475 0.2550 ;
        RECT 1.8600 0.1800 1.9425 0.2550 ;
        RECT 1.7850 0.1800 1.8600 0.3300 ;
        RECT 1.7325 0.7050 1.8375 0.8100 ;
        RECT 1.5000 0.2550 1.7850 0.3300 ;
        RECT 1.6875 0.4050 1.7775 0.6000 ;
        RECT 1.6200 0.7050 1.7325 0.7875 ;
        RECT 1.5975 0.4050 1.6875 0.5775 ;
        RECT 1.4700 0.6600 1.6200 0.7875 ;
        RECT 0.8400 0.4725 1.5225 0.5775 ;
        RECT 0.9150 0.2775 1.3950 0.3975 ;
        RECT 0.9150 0.6525 1.3950 0.7725 ;
        RECT 0.7650 0.3000 0.8400 0.7950 ;
        RECT 0.2550 0.3000 0.7650 0.3750 ;
        RECT 0.5775 0.7200 0.7650 0.7950 ;
        RECT 0.5250 0.4500 0.6900 0.6450 ;
        RECT 0.1575 0.1500 0.5850 0.2250 ;
        RECT 0.4725 0.7200 0.5775 0.8400 ;
        RECT 0.3975 0.4500 0.4500 0.6375 ;
        RECT 0.3075 0.4500 0.3975 0.7500 ;
        RECT 0.0525 0.1500 0.1575 0.2550 ;
        LAYER VIA1 ;
        RECT 1.5450 0.2550 1.6200 0.3300 ;
        RECT 1.5075 0.6750 1.5825 0.7500 ;
        RECT 0.5925 0.4950 0.6675 0.5700 ;
        LAYER M2 ;
        RECT 1.5675 0.2550 1.6650 0.3300 ;
        RECT 1.5675 0.6375 1.5975 0.7875 ;
        RECT 1.4925 0.1125 1.5675 0.7875 ;
        RECT 0.6825 0.1125 1.4925 0.1875 ;
        RECT 0.5775 0.1125 0.6825 0.6150 ;
    END
END MAOI22_0111


MACRO MAOI22_1000
    CLASS CORE ;
    FOREIGN MAOI22_1000 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.2600 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 0.7275 0.2625 0.8325 0.7725 ;
        RECT 0.2625 0.2625 0.7275 0.3375 ;
        VIA 0.7800 0.6825 VIA12_square ;
        VIA 0.7125 0.3000 VIA12_square ;
        END
    END ZN
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.4575 0.8625 0.6525 0.9375 ;
        RECT 0.3525 0.4800 0.4575 0.9375 ;
        RECT 0.0825 0.8625 0.3525 0.9375 ;
        VIA 0.4050 0.5625 VIA12_square ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1425 0.4500 0.2325 0.5700 ;
        RECT 0.0675 0.3675 0.1425 0.6825 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.1175 0.3675 1.1925 0.6825 ;
        RECT 1.0275 0.4350 1.1175 0.5550 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.9075 0.1125 1.0125 0.3225 ;
        RECT 0.4425 0.1125 0.9075 0.1875 ;
        VIA 0.9600 0.2400 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.2225 -0.0750 1.2600 0.0750 ;
        RECT 1.1175 -0.0750 1.2225 0.2475 ;
        RECT 0.5850 -0.0750 1.1175 0.0750 ;
        RECT 0.4650 -0.0750 0.5850 0.1800 ;
        RECT 0.1650 -0.0750 0.4650 0.0750 ;
        RECT 0.0450 -0.0750 0.1650 0.2475 ;
        RECT 0.0000 -0.0750 0.0450 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.5850 0.9750 1.2600 1.1250 ;
        RECT 0.4650 0.8700 0.5850 1.1250 ;
        RECT 0.0000 0.9750 0.4650 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.1250 0.1575 1.1850 0.2175 ;
        RECT 1.1250 0.8175 1.1850 0.8775 ;
        RECT 1.0275 0.4650 1.0875 0.5250 ;
        RECT 0.9150 0.6750 0.9750 0.7350 ;
        RECT 0.8100 0.4875 0.8700 0.5475 ;
        RECT 0.7050 0.1575 0.7650 0.2175 ;
        RECT 0.7050 0.8175 0.7650 0.8775 ;
        RECT 0.6000 0.4875 0.6600 0.5475 ;
        RECT 0.4950 0.1200 0.5550 0.1800 ;
        RECT 0.4950 0.8700 0.5550 0.9300 ;
        RECT 0.2850 0.1725 0.3450 0.2325 ;
        RECT 0.1725 0.4800 0.2325 0.5400 ;
        RECT 0.0750 0.1575 0.1350 0.2175 ;
        RECT 0.0750 0.8175 0.1350 0.8775 ;
        RECT 0.3825 0.4950 0.4425 0.5550 ;
        LAYER M1 ;
        RECT 1.1025 0.7950 1.2075 0.9000 ;
        RECT 0.7875 0.8250 1.1025 0.9000 ;
        RECT 0.9525 0.2025 1.0425 0.3600 ;
        RECT 0.8475 0.6450 1.0425 0.7500 ;
        RECT 0.8775 0.2025 0.9525 0.5700 ;
        RECT 0.7875 0.4650 0.8775 0.5700 ;
        RECT 0.6975 0.6450 0.8475 0.7200 ;
        RECT 0.6675 0.1500 0.8025 0.3900 ;
        RECT 0.6825 0.7950 0.7875 0.9000 ;
        RECT 0.5925 0.4650 0.6825 0.5700 ;
        RECT 0.5175 0.2550 0.5925 0.7950 ;
        RECT 0.3750 0.2550 0.5175 0.3300 ;
        RECT 0.3750 0.7200 0.5175 0.7950 ;
        RECT 0.3075 0.4050 0.4425 0.6450 ;
        RECT 0.2550 0.1500 0.3750 0.3300 ;
        RECT 0.3000 0.7200 0.3750 0.8700 ;
        RECT 0.1575 0.7950 0.3000 0.8700 ;
        RECT 0.0450 0.7950 0.1575 0.9000 ;
    END
END MAOI22_1000


MACRO MAOI22_1010
    CLASS CORE ;
    FOREIGN MAOI22_1010 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.2600 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 0.7875 0.6300 0.8550 0.7350 ;
        RECT 0.7050 0.2625 0.7875 0.7350 ;
        RECT 0.3150 0.2625 0.7050 0.3375 ;
        VIA 0.7800 0.6825 VIA12_square ;
        VIA 0.7425 0.3450 VIA12_square ;
        END
    END ZN
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.4575 0.7125 0.5325 0.7875 ;
        RECT 0.3675 0.4500 0.4575 0.7875 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.2100 0.4650 0.2925 0.8325 ;
        RECT 0.1875 0.4650 0.2100 0.5850 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.1175 0.3675 1.1925 0.6825 ;
        RECT 1.0275 0.4350 1.1175 0.5550 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.0125 0.1125 1.0950 0.1875 ;
        RECT 0.9075 0.1125 1.0125 0.3225 ;
        RECT 0.6300 0.1125 0.9075 0.1875 ;
        VIA 0.9600 0.2400 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.2225 -0.0750 1.2600 0.0750 ;
        RECT 1.1175 -0.0750 1.2225 0.2475 ;
        RECT 0.5850 -0.0750 1.1175 0.0750 ;
        RECT 0.4650 -0.0750 0.5850 0.1950 ;
        RECT 0.1650 -0.0750 0.4650 0.0750 ;
        RECT 0.0450 -0.0750 0.1650 0.2175 ;
        RECT 0.0000 -0.0750 0.0450 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.5850 0.9750 1.2600 1.1250 ;
        RECT 0.4650 0.8700 0.5850 1.1250 ;
        RECT 0.0000 0.9750 0.4650 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.1250 0.1575 1.1850 0.2175 ;
        RECT 1.1250 0.8175 1.1850 0.8775 ;
        RECT 1.0275 0.4650 1.0875 0.5250 ;
        RECT 0.9150 0.6750 0.9750 0.7350 ;
        RECT 0.8175 0.4950 0.8775 0.5550 ;
        RECT 0.7050 0.2400 0.7650 0.3000 ;
        RECT 0.7050 0.8175 0.7650 0.8775 ;
        RECT 0.5925 0.4950 0.6525 0.5550 ;
        RECT 0.4950 0.1275 0.5550 0.1875 ;
        RECT 0.4950 0.8700 0.5550 0.9300 ;
        RECT 0.3900 0.4800 0.4500 0.5400 ;
        RECT 0.2850 0.2775 0.3450 0.3375 ;
        RECT 0.1875 0.4950 0.2475 0.5550 ;
        RECT 0.0750 0.1575 0.1350 0.2175 ;
        RECT 0.0750 0.7800 0.1350 0.8400 ;
        LAYER M1 ;
        RECT 1.1025 0.7950 1.2075 0.9000 ;
        RECT 0.7875 0.8250 1.1025 0.9000 ;
        RECT 0.9525 0.2025 1.0425 0.3600 ;
        RECT 0.8475 0.6450 1.0425 0.7500 ;
        RECT 0.8775 0.2025 0.9525 0.5700 ;
        RECT 0.7875 0.4950 0.8775 0.5700 ;
        RECT 0.6525 0.6450 0.8475 0.7200 ;
        RECT 0.6825 0.1500 0.8025 0.4200 ;
        RECT 0.6825 0.7950 0.7875 0.9000 ;
        RECT 0.6075 0.4950 0.6825 0.5700 ;
        RECT 0.5325 0.2700 0.6075 0.5700 ;
        RECT 0.2925 0.2700 0.5325 0.3450 ;
        RECT 0.2250 0.2700 0.2925 0.3750 ;
        RECT 0.1125 0.3000 0.2250 0.3750 ;
        RECT 0.1125 0.7500 0.1350 0.8700 ;
        RECT 0.0375 0.3000 0.1125 0.8700 ;
    END
END MAOI22_1010


MACRO MOAI22_0011
    CLASS CORE ;
    FOREIGN MOAI22_0011 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.6800 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 0.9600 0.2625 1.0350 0.7875 ;
        RECT 0.4950 0.2625 0.9600 0.3375 ;
        RECT 0.8700 0.6825 0.9600 0.7875 ;
        VIA 0.9525 0.3000 VIA12_square ;
        VIA 0.9525 0.7350 VIA12_square ;
        END
    END ZN
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1425 0.4500 0.2325 0.5700 ;
        RECT 0.0675 0.3675 0.1425 0.6825 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.4575 0.7125 0.5325 0.7875 ;
        RECT 0.3525 0.4350 0.4575 0.7875 ;
        RECT 0.0675 0.7125 0.3525 0.7875 ;
        VIA 0.3975 0.5175 VIA12_square ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.1550 0.5625 1.6200 0.6375 ;
        VIA 1.4400 0.6000 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.1625 0.1125 1.2675 0.4200 ;
        RECT 0.6975 0.1125 1.1625 0.1875 ;
        VIA 1.2150 0.3375 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.6350 -0.0750 1.6800 0.0750 ;
        RECT 1.5150 -0.0750 1.6350 0.2175 ;
        RECT 1.2150 -0.0750 1.5150 0.0750 ;
        RECT 1.0950 -0.0750 1.2150 0.1800 ;
        RECT 0.7950 -0.0750 1.0950 0.0750 ;
        RECT 0.6750 -0.0750 0.7950 0.1800 ;
        RECT 0.1575 -0.0750 0.6750 0.0750 ;
        RECT 0.0525 -0.0750 0.1575 0.2400 ;
        RECT 0.0000 -0.0750 0.0525 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.2150 0.9750 1.6800 1.1250 ;
        RECT 1.0950 0.8625 1.2150 1.1250 ;
        RECT 0.8025 0.9750 1.0950 1.1250 ;
        RECT 0.6900 0.8400 0.8025 1.1250 ;
        RECT 0.0000 0.9750 0.6900 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.5450 0.1575 1.6050 0.2175 ;
        RECT 1.5450 0.8250 1.6050 0.8850 ;
        RECT 1.4325 0.4875 1.4925 0.5475 ;
        RECT 1.3350 0.2475 1.3950 0.3075 ;
        RECT 1.2300 0.4725 1.2900 0.5325 ;
        RECT 1.1250 0.1200 1.1850 0.1800 ;
        RECT 1.1250 0.8700 1.1850 0.9300 ;
        RECT 1.0200 0.4950 1.0800 0.5550 ;
        RECT 0.9150 0.2475 0.9750 0.3075 ;
        RECT 0.9150 0.6825 0.9750 0.7425 ;
        RECT 0.8100 0.4950 0.8700 0.5550 ;
        RECT 0.7050 0.1200 0.7650 0.1800 ;
        RECT 0.7050 0.8700 0.7650 0.9300 ;
        RECT 0.6000 0.4950 0.6600 0.5550 ;
        RECT 0.4950 0.2100 0.5550 0.2700 ;
        RECT 0.4950 0.8325 0.5550 0.8925 ;
        RECT 0.3900 0.4950 0.4500 0.5550 ;
        RECT 0.2850 0.6825 0.3450 0.7425 ;
        RECT 0.1725 0.4800 0.2325 0.5400 ;
        RECT 0.0750 0.1575 0.1350 0.2175 ;
        RECT 0.0750 0.8175 0.1350 0.8775 ;
        LAYER M1 ;
        RECT 1.5675 0.2925 1.6425 0.8925 ;
        RECT 1.4025 0.2925 1.5675 0.3675 ;
        RECT 1.3200 0.8175 1.5675 0.8925 ;
        RECT 1.3800 0.4425 1.4925 0.7425 ;
        RECT 1.3275 0.2025 1.4025 0.3675 ;
        RECT 1.2525 0.4425 1.2975 0.5775 ;
        RECT 1.1775 0.2550 1.2525 0.5775 ;
        RECT 1.1325 0.2550 1.1775 0.3600 ;
        RECT 1.0200 0.6525 1.1175 0.7800 ;
        RECT 0.8400 0.4725 1.1025 0.5775 ;
        RECT 1.0200 0.2475 1.0575 0.3975 ;
        RECT 0.9150 0.1500 1.0200 0.3975 ;
        RECT 0.9150 0.6525 1.0200 0.9000 ;
        RECT 0.7650 0.2550 0.8400 0.7500 ;
        RECT 0.5625 0.2550 0.7650 0.3300 ;
        RECT 0.2550 0.6750 0.7650 0.7500 ;
        RECT 0.5250 0.4050 0.6900 0.6000 ;
        RECT 0.1575 0.8250 0.5850 0.9000 ;
        RECT 0.4875 0.1725 0.5625 0.3300 ;
        RECT 0.3975 0.4050 0.4500 0.6000 ;
        RECT 0.3075 0.2850 0.3975 0.6000 ;
        RECT 0.0525 0.7950 0.1575 0.9000 ;
        LAYER VIA1 ;
        RECT 1.3650 0.8175 1.4400 0.8925 ;
        RECT 0.5925 0.4800 0.6675 0.5550 ;
        LAYER M2 ;
        RECT 1.2975 0.8175 1.4850 0.9375 ;
        RECT 0.7725 0.8625 1.2975 0.9375 ;
        RECT 0.6975 0.4650 0.7725 0.9375 ;
        RECT 0.5475 0.4650 0.6975 0.5700 ;
    END
END MOAI22_0011


MACRO MOAI22_0100
    CLASS CORE ;
    FOREIGN MOAI22_0100 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.0900 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 1.7400 0.2625 2.0550 0.7800 ;
        VIA 1.8975 0.3450 VIA12_slot ;
        VIA 1.8975 0.6975 VIA12_slot ;
        END
    END ZN
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 5.9475 0.4050 6.0225 0.6900 ;
        RECT 5.8575 0.4050 5.9475 0.5700 ;
        RECT 4.7700 0.4650 5.8575 0.5700 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 4.0950 0.4125 4.4550 0.4875 ;
        RECT 3.9900 0.4125 4.0950 0.6375 ;
        VIA 4.0425 0.5250 VIA12_square ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.2775 0.4650 1.2825 0.5850 ;
        RECT 0.1425 0.4650 0.2775 0.6450 ;
        RECT 0.0675 0.3675 0.1425 0.6450 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.4850 0.4500 1.5900 0.6375 ;
        RECT 1.0650 0.5325 1.4850 0.6375 ;
        VIA 1.5375 0.5325 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 5.8350 -0.0750 6.0900 0.0750 ;
        RECT 5.7150 -0.0750 5.8350 0.1800 ;
        RECT 5.4150 -0.0750 5.7150 0.0750 ;
        RECT 5.2950 -0.0750 5.4150 0.1800 ;
        RECT 4.9950 -0.0750 5.2950 0.0750 ;
        RECT 4.8750 -0.0750 4.9950 0.1800 ;
        RECT 3.3075 -0.0750 4.8750 0.0750 ;
        RECT 3.2025 -0.0750 3.3075 0.2250 ;
        RECT 2.8875 -0.0750 3.2025 0.0750 ;
        RECT 2.7825 -0.0750 2.8875 0.2250 ;
        RECT 2.4675 -0.0750 2.7825 0.0750 ;
        RECT 2.3625 -0.0750 2.4675 0.2250 ;
        RECT 0.0000 -0.0750 2.3625 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 6.0375 0.9750 6.0900 1.1250 ;
        RECT 5.9325 0.8100 6.0375 1.1250 ;
        RECT 5.6250 0.9750 5.9325 1.1250 ;
        RECT 5.5050 0.8325 5.6250 1.1250 ;
        RECT 5.2050 0.9750 5.5050 1.1250 ;
        RECT 5.0850 0.8325 5.2050 1.1250 ;
        RECT 4.7850 0.9750 5.0850 1.1250 ;
        RECT 4.6650 0.8325 4.7850 1.1250 ;
        RECT 4.3650 0.9750 4.6650 1.1250 ;
        RECT 4.2450 0.8700 4.3650 1.1250 ;
        RECT 3.9450 0.9750 4.2450 1.1250 ;
        RECT 3.8250 0.8325 3.9450 1.1250 ;
        RECT 3.3075 0.9750 3.8250 1.1250 ;
        RECT 3.2025 0.8250 3.3075 1.1250 ;
        RECT 2.8875 0.9750 3.2025 1.1250 ;
        RECT 2.7825 0.8250 2.8875 1.1250 ;
        RECT 1.2150 0.9750 2.7825 1.1250 ;
        RECT 1.0950 0.8700 1.2150 1.1250 ;
        RECT 0.7950 0.9750 1.0950 1.1250 ;
        RECT 0.6750 0.8700 0.7950 1.1250 ;
        RECT 0.3750 0.9750 0.6750 1.1250 ;
        RECT 0.2550 0.8700 0.3750 1.1250 ;
        RECT 0.0000 0.9750 0.2550 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 5.9550 0.2400 6.0150 0.3000 ;
        RECT 5.9550 0.8325 6.0150 0.8925 ;
        RECT 5.8500 0.4950 5.9100 0.5550 ;
        RECT 5.7450 0.1200 5.8050 0.1800 ;
        RECT 5.7450 0.7500 5.8050 0.8100 ;
        RECT 5.6400 0.4950 5.7000 0.5550 ;
        RECT 5.5350 0.2850 5.5950 0.3450 ;
        RECT 5.5350 0.8325 5.5950 0.8925 ;
        RECT 5.4300 0.4950 5.4900 0.5550 ;
        RECT 5.3250 0.1200 5.3850 0.1800 ;
        RECT 5.3250 0.7500 5.3850 0.8100 ;
        RECT 5.2200 0.4950 5.2800 0.5550 ;
        RECT 5.1150 0.3075 5.1750 0.3675 ;
        RECT 5.1150 0.8325 5.1750 0.8925 ;
        RECT 5.0100 0.4950 5.0700 0.5550 ;
        RECT 4.9050 0.1200 4.9650 0.1800 ;
        RECT 4.8000 0.4950 4.8600 0.5550 ;
        RECT 4.6950 0.2250 4.7550 0.2850 ;
        RECT 4.6950 0.8325 4.7550 0.8925 ;
        RECT 4.5900 0.4950 4.6500 0.5550 ;
        RECT 4.4850 0.3075 4.5450 0.3675 ;
        RECT 4.4850 0.7500 4.5450 0.8100 ;
        RECT 4.3800 0.4950 4.4400 0.5550 ;
        RECT 4.2750 0.1575 4.3350 0.2175 ;
        RECT 4.2750 0.8700 4.3350 0.9300 ;
        RECT 4.1700 0.4950 4.2300 0.5550 ;
        RECT 4.0650 0.3075 4.1250 0.3675 ;
        RECT 4.0650 0.7275 4.1250 0.7875 ;
        RECT 3.9600 0.4950 4.0200 0.5550 ;
        RECT 3.8550 0.1575 3.9150 0.2175 ;
        RECT 3.8550 0.8325 3.9150 0.8925 ;
        RECT 3.7500 0.4950 3.8100 0.5550 ;
        RECT 3.6450 0.3075 3.7050 0.3675 ;
        RECT 3.4350 0.2775 3.4950 0.3375 ;
        RECT 3.4350 0.7275 3.4950 0.7875 ;
        RECT 3.3300 0.4950 3.3900 0.5550 ;
        RECT 3.2250 0.1425 3.2850 0.2025 ;
        RECT 3.2250 0.8475 3.2850 0.9075 ;
        RECT 3.1200 0.4950 3.1800 0.5550 ;
        RECT 3.0150 0.3075 3.0750 0.3675 ;
        RECT 3.0150 0.6900 3.0750 0.7500 ;
        RECT 2.9100 0.4950 2.9700 0.5550 ;
        RECT 2.8050 0.1425 2.8650 0.2025 ;
        RECT 2.8050 0.8475 2.8650 0.9075 ;
        RECT 2.7000 0.4950 2.7600 0.5550 ;
        RECT 2.5950 0.3075 2.6550 0.3675 ;
        RECT 2.5950 0.6900 2.6550 0.7500 ;
        RECT 2.4900 0.4950 2.5500 0.5550 ;
        RECT 2.3850 0.1425 2.4450 0.2025 ;
        RECT 2.2800 0.4950 2.3400 0.5550 ;
        RECT 2.1750 0.2400 2.2350 0.3000 ;
        RECT 2.1750 0.8325 2.2350 0.8925 ;
        RECT 2.0625 0.4950 2.1225 0.5550 ;
        RECT 1.9650 0.3075 2.0250 0.3675 ;
        RECT 1.9650 0.6900 2.0250 0.7500 ;
        RECT 1.8600 0.4950 1.9200 0.5550 ;
        RECT 1.7550 0.1575 1.8150 0.2175 ;
        RECT 1.7550 0.8325 1.8150 0.8925 ;
        RECT 1.6500 0.4950 1.7100 0.5550 ;
        RECT 1.5450 0.3075 1.6050 0.3675 ;
        RECT 1.5450 0.6900 1.6050 0.7500 ;
        RECT 1.4400 0.4950 1.5000 0.5550 ;
        RECT 1.3350 0.1575 1.3950 0.2175 ;
        RECT 1.3350 0.7575 1.3950 0.8175 ;
        RECT 1.2225 0.4950 1.2825 0.5550 ;
        RECT 1.1250 0.3075 1.1850 0.3675 ;
        RECT 1.1250 0.8700 1.1850 0.9300 ;
        RECT 1.0200 0.4950 1.0800 0.5550 ;
        RECT 0.9150 0.1575 0.9750 0.2175 ;
        RECT 0.9150 0.7275 0.9750 0.7875 ;
        RECT 0.8100 0.4950 0.8700 0.5550 ;
        RECT 0.7050 0.8700 0.7650 0.9300 ;
        RECT 0.6000 0.4950 0.6600 0.5550 ;
        RECT 0.4950 0.1575 0.5550 0.2175 ;
        RECT 0.4950 0.7275 0.5550 0.7875 ;
        RECT 0.3900 0.4950 0.4500 0.5550 ;
        RECT 0.2850 0.3225 0.3450 0.3825 ;
        RECT 0.2850 0.8700 0.3450 0.9300 ;
        RECT 0.1800 0.4950 0.2400 0.5550 ;
        RECT 0.0750 0.1725 0.1350 0.2325 ;
        RECT 0.0750 0.7575 0.1350 0.8175 ;
        LAYER M1 ;
        RECT 5.9475 0.2100 6.0225 0.3300 ;
        RECT 5.6025 0.2550 5.9475 0.3300 ;
        RECT 5.7375 0.6450 5.8125 0.8475 ;
        RECT 5.3925 0.6450 5.7375 0.7575 ;
        RECT 5.5275 0.2550 5.6025 0.3750 ;
        RECT 4.7625 0.3000 5.5275 0.3750 ;
        RECT 5.3175 0.6450 5.3925 0.8475 ;
        RECT 4.5525 0.6450 5.3175 0.7575 ;
        RECT 4.6875 0.1500 4.7625 0.3750 ;
        RECT 3.8100 0.1500 4.6875 0.2250 ;
        RECT 3.7200 0.4650 4.6800 0.5700 ;
        RECT 3.6450 0.3000 4.5825 0.3750 ;
        RECT 4.4775 0.6450 4.5525 0.8475 ;
        RECT 4.1325 0.6450 4.4775 0.7575 ;
        RECT 4.0575 0.6450 4.1325 0.8475 ;
        RECT 3.6450 0.6450 4.0575 0.7500 ;
        RECT 3.5700 0.3000 3.6450 0.7500 ;
        RECT 2.2425 0.4650 3.5700 0.5700 ;
        RECT 3.4200 0.2400 3.4950 0.3750 ;
        RECT 3.4200 0.6450 3.4950 0.8250 ;
        RECT 2.2425 0.3000 3.4200 0.3750 ;
        RECT 1.5150 0.6450 3.4200 0.7500 ;
        RECT 1.4025 0.8250 2.2800 0.9000 ;
        RECT 2.1675 0.1500 2.2425 0.3750 ;
        RECT 0.1575 0.1500 2.1675 0.2250 ;
        RECT 1.3950 0.4650 2.1525 0.5700 ;
        RECT 0.2475 0.3000 2.0625 0.3900 ;
        RECT 1.3275 0.7200 1.4025 0.9000 ;
        RECT 0.1425 0.7200 1.3275 0.7950 ;
        RECT 0.0525 0.1500 0.1575 0.2550 ;
        RECT 0.0675 0.7200 0.1425 0.8475 ;
    END
END MOAI22_0100


MACRO MOAI22_0111
    CLASS CORE ;
    FOREIGN MOAI22_0111 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.1000 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 0.9975 0.2700 1.3125 0.7800 ;
        VIA 1.1550 0.3525 VIA12_slot ;
        VIA 1.1550 0.6975 VIA12_slot ;
        END
    END ZN
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1425 0.4500 0.2325 0.5700 ;
        RECT 0.0675 0.3675 0.1425 0.6825 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.4575 0.7125 0.6675 0.7875 ;
        RECT 0.3525 0.4350 0.4575 0.7875 ;
        RECT 0.1275 0.7125 0.3525 0.7875 ;
        VIA 0.3975 0.5175 VIA12_square ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.9575 0.3675 2.0325 0.6825 ;
        RECT 1.8600 0.4500 1.9575 0.5700 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.7475 0.8625 2.0250 0.9375 ;
        RECT 1.6725 0.4125 1.7475 0.9375 ;
        RECT 1.6425 0.4125 1.6725 0.5625 ;
        RECT 1.4700 0.8625 1.6725 0.9375 ;
        VIA 1.6950 0.4875 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 2.0475 -0.0750 2.1000 0.0750 ;
        RECT 1.9425 -0.0750 2.0475 0.2400 ;
        RECT 1.6350 -0.0750 1.9425 0.0750 ;
        RECT 1.5150 -0.0750 1.6350 0.1800 ;
        RECT 1.2150 -0.0750 1.5150 0.0750 ;
        RECT 1.0950 -0.0750 1.2150 0.2025 ;
        RECT 0.7950 -0.0750 1.0950 0.0750 ;
        RECT 0.6750 -0.0750 0.7950 0.1800 ;
        RECT 0.1575 -0.0750 0.6750 0.0750 ;
        RECT 0.0525 -0.0750 0.1575 0.2400 ;
        RECT 0.0000 -0.0750 0.0525 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.6350 0.9750 2.1000 1.1250 ;
        RECT 1.5150 0.8625 1.6350 1.1250 ;
        RECT 1.2150 0.9750 1.5150 1.1250 ;
        RECT 1.0950 0.8475 1.2150 1.1250 ;
        RECT 0.8025 0.9750 1.0950 1.1250 ;
        RECT 0.6900 0.8400 0.8025 1.1250 ;
        RECT 0.0000 0.9750 0.6900 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.9650 0.1575 2.0250 0.2175 ;
        RECT 1.9650 0.8175 2.0250 0.8775 ;
        RECT 1.8600 0.4800 1.9200 0.5400 ;
        RECT 1.7550 0.1725 1.8150 0.2325 ;
        RECT 1.6500 0.4800 1.7100 0.5400 ;
        RECT 1.5450 0.1200 1.6050 0.1800 ;
        RECT 1.5450 0.8700 1.6050 0.9300 ;
        RECT 1.4400 0.4950 1.5000 0.5550 ;
        RECT 1.3350 0.3075 1.3950 0.3675 ;
        RECT 1.3350 0.6825 1.3950 0.7425 ;
        RECT 1.2300 0.4950 1.2900 0.5550 ;
        RECT 1.1250 0.1350 1.1850 0.1950 ;
        RECT 1.1250 0.8550 1.1850 0.9150 ;
        RECT 1.0200 0.4950 1.0800 0.5550 ;
        RECT 0.9150 0.3075 0.9750 0.3675 ;
        RECT 0.9150 0.6825 0.9750 0.7425 ;
        RECT 0.8100 0.4950 0.8700 0.5550 ;
        RECT 0.7050 0.1200 0.7650 0.1800 ;
        RECT 0.7050 0.8700 0.7650 0.9300 ;
        RECT 0.6000 0.4950 0.6600 0.5550 ;
        RECT 0.4950 0.2100 0.5550 0.2700 ;
        RECT 0.4950 0.8325 0.5550 0.8925 ;
        RECT 0.3900 0.4950 0.4500 0.5550 ;
        RECT 0.2850 0.6825 0.3450 0.7425 ;
        RECT 0.1725 0.4800 0.2325 0.5400 ;
        RECT 0.0750 0.1575 0.1350 0.2175 ;
        RECT 0.0750 0.8175 0.1350 0.8775 ;
        LAYER M1 ;
        RECT 1.8450 0.7950 2.0475 0.9000 ;
        RECT 1.7625 0.7050 1.8450 0.9000 ;
        RECT 1.8075 0.1500 1.8375 0.2550 ;
        RECT 1.7325 0.1500 1.8075 0.3300 ;
        RECT 1.6875 0.4050 1.7775 0.6000 ;
        RECT 1.6200 0.7050 1.7625 0.7875 ;
        RECT 1.5000 0.2550 1.7325 0.3300 ;
        RECT 1.5975 0.4050 1.6875 0.5775 ;
        RECT 1.4700 0.6600 1.6200 0.7875 ;
        RECT 0.8400 0.4725 1.5225 0.5775 ;
        RECT 0.9150 0.2775 1.3950 0.3975 ;
        RECT 0.9150 0.6525 1.3950 0.7725 ;
        RECT 0.7650 0.2550 0.8400 0.7500 ;
        RECT 0.5625 0.2550 0.7650 0.3300 ;
        RECT 0.2550 0.6750 0.7650 0.7500 ;
        RECT 0.5250 0.4050 0.6900 0.6000 ;
        RECT 0.1575 0.8250 0.5850 0.9000 ;
        RECT 0.4875 0.1725 0.5625 0.3300 ;
        RECT 0.3975 0.4050 0.4500 0.6000 ;
        RECT 0.3075 0.2850 0.3975 0.6000 ;
        RECT 0.0525 0.7950 0.1575 0.9000 ;
        LAYER VIA1 ;
        RECT 1.5450 0.2550 1.6200 0.3300 ;
        RECT 1.5075 0.6750 1.5825 0.7500 ;
        RECT 0.5925 0.4500 0.6675 0.5250 ;
        LAYER M2 ;
        RECT 1.5675 0.2550 1.6650 0.3300 ;
        RECT 1.5675 0.6375 1.5975 0.7875 ;
        RECT 1.4925 0.1125 1.5675 0.7875 ;
        RECT 0.6825 0.1125 1.4925 0.1875 ;
        RECT 0.5775 0.1125 0.6825 0.5700 ;
    END
END MOAI22_0111


MACRO MOAI22_1000
    CLASS CORE ;
    FOREIGN MOAI22_1000 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.2600 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 0.8025 0.1125 0.8775 0.7875 ;
        RECT 0.3075 0.1125 0.8025 0.1875 ;
        RECT 0.6225 0.7125 0.8025 0.7875 ;
        VIA 0.8400 0.3675 VIA12_square ;
        VIA 0.7050 0.7500 VIA12_square ;
        END
    END ZN
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.4275 0.2625 0.6075 0.3375 ;
        RECT 0.3525 0.2625 0.4275 0.5700 ;
        RECT 0.0675 0.2625 0.3525 0.3375 ;
        VIA 0.3900 0.4875 VIA12_square ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1575 0.4500 0.2325 0.5700 ;
        RECT 0.0525 0.3675 0.1575 0.6825 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.1175 0.3675 1.2075 0.6825 ;
        RECT 0.9975 0.4950 1.1175 0.6000 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.0575 0.8625 1.1925 0.9375 ;
        RECT 0.9525 0.7125 1.0575 0.9375 ;
        RECT 0.6525 0.8625 0.9525 0.9375 ;
        VIA 1.0050 0.7875 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.5850 -0.0750 1.2600 0.0750 ;
        RECT 0.4650 -0.0750 0.5850 0.1800 ;
        RECT 0.0000 -0.0750 0.4650 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.2225 0.9750 1.2600 1.1250 ;
        RECT 1.1175 0.8025 1.2225 1.1250 ;
        RECT 0.5850 0.9750 1.1175 1.1250 ;
        RECT 0.4650 0.8700 0.5850 1.1250 ;
        RECT 0.1575 0.9750 0.4650 1.1250 ;
        RECT 0.0525 0.7950 0.1575 1.1250 ;
        RECT 0.0000 0.9750 0.0525 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.1250 0.1650 1.1850 0.2250 ;
        RECT 1.1250 0.8325 1.1850 0.8925 ;
        RECT 1.0275 0.4950 1.0875 0.5550 ;
        RECT 0.9150 0.3000 0.9750 0.3600 ;
        RECT 0.8175 0.4950 0.8775 0.5550 ;
        RECT 0.7050 0.1575 0.7650 0.2175 ;
        RECT 0.7050 0.8325 0.7650 0.8925 ;
        RECT 0.5925 0.4875 0.6525 0.5475 ;
        RECT 0.4950 0.1200 0.5550 0.1800 ;
        RECT 0.4950 0.8700 0.5550 0.9300 ;
        RECT 0.3825 0.4800 0.4425 0.5400 ;
        RECT 0.2850 0.7950 0.3450 0.8550 ;
        RECT 0.1725 0.4800 0.2325 0.5400 ;
        RECT 0.0750 0.1575 0.1350 0.2175 ;
        RECT 0.0750 0.8250 0.1350 0.8850 ;
        LAYER M1 ;
        RECT 1.1100 0.1500 1.2150 0.2550 ;
        RECT 0.7725 0.1500 1.1100 0.2250 ;
        RECT 0.8325 0.3000 1.0425 0.4200 ;
        RECT 0.9675 0.6750 1.0425 0.8700 ;
        RECT 0.9225 0.6750 0.9675 0.7500 ;
        RECT 0.8475 0.4950 0.9225 0.7500 ;
        RECT 0.7725 0.8250 0.8625 0.9000 ;
        RECT 0.7875 0.4950 0.8475 0.5700 ;
        RECT 0.7350 0.3300 0.8325 0.4200 ;
        RECT 0.6675 0.1500 0.7725 0.2550 ;
        RECT 0.6675 0.6450 0.7725 0.9000 ;
        RECT 0.5925 0.4650 0.6750 0.5700 ;
        RECT 0.5175 0.2550 0.5925 0.7950 ;
        RECT 0.3900 0.2550 0.5175 0.3300 ;
        RECT 0.3600 0.7200 0.5175 0.7950 ;
        RECT 0.3075 0.4050 0.4425 0.6450 ;
        RECT 0.3150 0.1875 0.3900 0.3300 ;
        RECT 0.2550 0.7200 0.3600 0.8850 ;
        RECT 0.1650 0.1875 0.3150 0.2925 ;
        RECT 0.0450 0.1500 0.1650 0.2925 ;
    END
END MOAI22_1000


MACRO MOAI22_1010
    CLASS CORE ;
    FOREIGN MOAI22_1010 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.2600 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 0.8175 0.2850 0.8475 0.3900 ;
        RECT 0.7425 0.2850 0.8175 0.7875 ;
        RECT 0.3525 0.7125 0.7425 0.7875 ;
        VIA 0.7800 0.3675 VIA12_square ;
        VIA 0.7350 0.7500 VIA12_square ;
        END
    END ZN
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.0675 0.4125 0.5325 0.4875 ;
        VIA 0.4050 0.4500 VIA12_square ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.0675 0.2625 0.5325 0.3375 ;
        VIA 0.2475 0.3000 VIA12_square ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.1175 0.3675 1.2075 0.6825 ;
        RECT 1.0275 0.4650 1.1175 0.5850 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.9975 0.8625 1.0950 0.9375 ;
        RECT 0.8925 0.7125 0.9975 0.9375 ;
        RECT 0.5550 0.8625 0.8925 0.9375 ;
        VIA 0.9450 0.7875 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.5850 -0.0750 1.2600 0.0750 ;
        RECT 0.4650 -0.0750 0.5850 0.1875 ;
        RECT 0.0000 -0.0750 0.4650 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.2225 0.9750 1.2600 1.1250 ;
        RECT 1.1175 0.8025 1.2225 1.1250 ;
        RECT 0.5850 0.9750 1.1175 1.1250 ;
        RECT 0.4650 0.8700 0.5850 1.1250 ;
        RECT 0.1650 0.9750 0.4650 1.1250 ;
        RECT 0.0450 0.8325 0.1650 1.1250 ;
        RECT 0.0000 0.9750 0.0450 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.1250 0.1650 1.1850 0.2250 ;
        RECT 1.1250 0.8325 1.1850 0.8925 ;
        RECT 1.0275 0.4950 1.0875 0.5550 ;
        RECT 0.9150 0.3000 0.9750 0.3600 ;
        RECT 0.8175 0.4950 0.8775 0.5550 ;
        RECT 0.7050 0.1575 0.7650 0.2175 ;
        RECT 0.7050 0.7500 0.7650 0.8100 ;
        RECT 0.5925 0.4950 0.6525 0.5550 ;
        RECT 0.4950 0.1275 0.5550 0.1875 ;
        RECT 0.4950 0.8700 0.5550 0.9300 ;
        RECT 0.3825 0.4800 0.4425 0.5400 ;
        RECT 0.2850 0.6900 0.3450 0.7500 ;
        RECT 0.1875 0.4800 0.2475 0.5400 ;
        RECT 0.0750 0.2100 0.1350 0.2700 ;
        RECT 0.0750 0.8325 0.1350 0.8925 ;
        LAYER M1 ;
        RECT 1.1100 0.1500 1.2150 0.2550 ;
        RECT 0.7800 0.1500 1.1100 0.2250 ;
        RECT 0.9150 0.3000 1.0050 0.3900 ;
        RECT 0.9525 0.7125 0.9975 0.8625 ;
        RECT 0.8775 0.4800 0.9525 0.8625 ;
        RECT 0.8400 0.3000 0.9150 0.4050 ;
        RECT 0.7875 0.4800 0.8775 0.5550 ;
        RECT 0.6300 0.3300 0.8400 0.4050 ;
        RECT 0.6750 0.6300 0.7950 0.9000 ;
        RECT 0.6750 0.1500 0.7800 0.2550 ;
        RECT 0.6000 0.4800 0.6825 0.5550 ;
        RECT 0.5250 0.4800 0.6000 0.7575 ;
        RECT 0.4500 0.2625 0.5250 0.3375 ;
        RECT 0.1125 0.6825 0.5250 0.7575 ;
        RECT 0.3600 0.2625 0.4500 0.5700 ;
        RECT 0.2100 0.1800 0.2850 0.5700 ;
        RECT 0.1875 0.3900 0.2100 0.5700 ;
        RECT 0.1125 0.1800 0.1350 0.3000 ;
        RECT 0.0375 0.1800 0.1125 0.7575 ;
    END
END MOAI22_1010


MACRO MUX2N_0011
    CLASS CORE ;
    FOREIGN MUX2N_0011 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.3100 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 1.9425 0.7725 2.0475 0.9375 ;
        RECT 1.3950 0.8625 1.9425 0.9375 ;
        RECT 1.3200 0.1125 1.3950 0.9375 ;
        RECT 0.7950 0.1125 1.3200 0.1875 ;
        RECT 0.7950 0.8625 1.3200 0.9375 ;
        RECT 0.6900 0.1125 0.7950 0.2775 ;
        RECT 0.6900 0.7725 0.7950 0.9375 ;
        VIA 1.9950 0.8475 VIA12_square ;
        VIA 1.3575 0.8475 VIA12_square ;
        VIA 1.3575 0.2025 VIA12_square ;
        VIA 0.7425 0.2025 VIA12_square ;
        VIA 0.7425 0.8475 VIA12_square ;
        END
    END ZN
    PIN S
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 2.0400 0.3150 2.1225 0.4350 ;
        RECT 1.7025 0.3150 2.0400 0.3900 ;
        RECT 1.6500 0.3150 1.7025 0.4050 ;
        RECT 1.3350 0.3300 1.6500 0.4050 ;
        RECT 1.2600 0.3300 1.3350 0.5700 ;
        RECT 0.8775 0.4950 1.2600 0.5700 ;
        RECT 0.8025 0.4950 0.8775 0.7200 ;
        RECT 0.3525 0.6450 0.8025 0.7200 ;
        RECT 0.2775 0.6450 0.3525 0.8325 ;
        RECT 0.2400 0.6450 0.2775 0.7200 ;
        RECT 0.0675 0.5175 0.2400 0.7200 ;
        END
    END S
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.9050 0.5625 2.2200 0.6375 ;
        RECT 1.8300 0.4125 1.9050 0.6375 ;
        RECT 1.5150 0.4125 1.8300 0.4875 ;
        VIA 1.8675 0.5175 VIA12_square ;
        END
    END I1
    PIN I0
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.5850 0.4125 1.0500 0.4875 ;
        RECT 0.4800 0.4125 0.5850 0.6075 ;
        VIA 0.5325 0.5250 VIA12_square ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.8375 -0.0750 2.3100 0.0750 ;
        RECT 1.7325 -0.0750 1.8375 0.2400 ;
        RECT 0.9975 -0.0750 1.7325 0.0750 ;
        RECT 0.8925 -0.0750 0.9975 0.2400 ;
        RECT 0.1575 -0.0750 0.8925 0.0750 ;
        RECT 0.0525 -0.0750 0.1575 0.2400 ;
        RECT 0.0000 -0.0750 0.0525 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.8375 0.9750 2.3100 1.1250 ;
        RECT 1.7325 0.8100 1.8375 1.1250 ;
        RECT 0.9975 0.9750 1.7325 1.1250 ;
        RECT 0.8925 0.8100 0.9975 1.1250 ;
        RECT 0.1575 0.9750 0.8925 1.1250 ;
        RECT 0.0525 0.8100 0.1575 1.1250 ;
        RECT 0.0000 0.9750 0.0525 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 2.1750 0.1575 2.2350 0.2175 ;
        RECT 2.1750 0.8175 2.2350 0.8775 ;
        RECT 2.0625 0.3450 2.1225 0.4050 ;
        RECT 2.0625 0.5850 2.1225 0.6450 ;
        RECT 1.8525 0.4875 1.9125 0.5475 ;
        RECT 1.7550 0.1575 1.8150 0.2175 ;
        RECT 1.7550 0.8325 1.8150 0.8925 ;
        RECT 1.6575 0.4950 1.7175 0.5550 ;
        RECT 1.4400 0.3450 1.5000 0.4050 ;
        RECT 1.4325 0.5850 1.4925 0.6450 ;
        RECT 1.3350 0.1725 1.3950 0.2325 ;
        RECT 1.3350 0.8175 1.3950 0.8775 ;
        RECT 1.1250 0.2025 1.1850 0.2625 ;
        RECT 1.1250 0.7425 1.1850 0.8025 ;
        RECT 1.0200 0.5025 1.0800 0.5625 ;
        RECT 0.9150 0.1575 0.9750 0.2175 ;
        RECT 0.9150 0.8325 0.9750 0.8925 ;
        RECT 0.8100 0.3450 0.8700 0.4050 ;
        RECT 0.8100 0.5850 0.8700 0.6450 ;
        RECT 0.6000 0.4950 0.6600 0.5550 ;
        RECT 0.4950 0.1725 0.5550 0.2325 ;
        RECT 0.4950 0.8175 0.5550 0.8775 ;
        RECT 0.3900 0.4950 0.4500 0.5550 ;
        RECT 0.1800 0.3450 0.2400 0.4050 ;
        RECT 0.1800 0.5850 0.2400 0.6450 ;
        RECT 0.0750 0.1575 0.1350 0.2175 ;
        RECT 0.0750 0.8325 0.1350 0.8925 ;
        LAYER M1 ;
        RECT 2.1975 0.1500 2.2725 0.9000 ;
        RECT 2.1375 0.1500 2.1975 0.2250 ;
        RECT 1.9200 0.7950 2.1975 0.9000 ;
        RECT 2.0475 0.5550 2.1225 0.7200 ;
        RECT 1.4925 0.6450 2.0475 0.7200 ;
        RECT 1.7700 0.4650 1.9425 0.5700 ;
        RECT 1.5975 0.4800 1.7700 0.5700 ;
        RECT 1.2675 0.7950 1.6575 0.9000 ;
        RECT 1.2600 0.1500 1.5600 0.2550 ;
        RECT 1.4175 0.5550 1.4925 0.7200 ;
        RECT 1.1850 0.6450 1.4175 0.7200 ;
        RECT 1.0800 0.1725 1.1850 0.4050 ;
        RECT 1.0800 0.6450 1.1850 0.8475 ;
        RECT 0.1500 0.3300 1.0800 0.4050 ;
        RECT 0.4725 0.1500 0.8175 0.2550 ;
        RECT 0.4725 0.7950 0.8175 0.9000 ;
        RECT 0.3450 0.4800 0.6975 0.5700 ;
        LAYER VIA1 ;
        RECT 1.1550 0.6450 1.2300 0.7200 ;
        RECT 1.0950 0.2625 1.1700 0.3375 ;
        LAYER M2 ;
        RECT 1.1700 0.2625 1.2450 0.7575 ;
        RECT 1.0200 0.2625 1.1700 0.3375 ;
        RECT 1.1400 0.6075 1.1700 0.7575 ;
    END
END MUX2N_0011


MACRO MUX2N_0111
    CLASS CORE ;
    FOREIGN MUX2N_0111 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.5200 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 1.8375 0.2850 2.1525 0.7275 ;
        VIA 1.9950 0.3450 VIA12_slot ;
        VIA 1.9950 0.6675 VIA12_slot ;
        END
    END ZN
    PIN S
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.6975 0.5625 1.1700 0.6375 ;
        RECT 0.5925 0.4725 0.6975 0.6375 ;
        VIA 0.6450 0.5475 VIA12_square ;
        END
    END S
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.9150 0.4125 1.3800 0.4875 ;
        VIA 1.0275 0.4500 VIA12_square ;
        END
    END I1
    PIN I0
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.4500 0.2625 0.9150 0.3375 ;
        VIA 0.5625 0.3000 VIA12_square ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 2.4525 -0.0750 2.5200 0.0750 ;
        RECT 2.3775 -0.0750 2.4525 0.3150 ;
        RECT 2.0550 -0.0750 2.3775 0.0750 ;
        RECT 1.9350 -0.0750 2.0550 0.1950 ;
        RECT 1.6350 -0.0750 1.9350 0.0750 ;
        RECT 1.5150 -0.0750 1.6350 0.1875 ;
        RECT 1.2150 -0.0750 1.5150 0.0750 ;
        RECT 1.0950 -0.0750 1.2150 0.1800 ;
        RECT 0.3750 -0.0750 1.0950 0.0750 ;
        RECT 0.2550 -0.0750 0.3750 0.2100 ;
        RECT 0.0000 -0.0750 0.2550 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 2.4525 0.9750 2.5200 1.1250 ;
        RECT 2.3775 0.6375 2.4525 1.1250 ;
        RECT 2.0325 0.9750 2.3775 1.1250 ;
        RECT 1.9575 0.8175 2.0325 1.1250 ;
        RECT 1.6350 0.9750 1.9575 1.1250 ;
        RECT 1.5150 0.8175 1.6350 1.1250 ;
        RECT 1.2225 0.9750 1.5150 1.1250 ;
        RECT 1.1175 0.8400 1.2225 1.1250 ;
        RECT 0.3750 0.9750 1.1175 1.1250 ;
        RECT 0.2550 0.8550 0.3750 1.1250 ;
        RECT 0.0000 0.9750 0.2550 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 2.3850 0.2250 2.4450 0.2850 ;
        RECT 2.3850 0.6675 2.4450 0.7275 ;
        RECT 2.3850 0.8325 2.4450 0.8925 ;
        RECT 2.2800 0.4650 2.3400 0.5250 ;
        RECT 2.1750 0.2250 2.2350 0.2850 ;
        RECT 2.1750 0.7200 2.2350 0.7800 ;
        RECT 2.0700 0.4650 2.1300 0.5250 ;
        RECT 1.9650 0.1275 2.0250 0.1875 ;
        RECT 1.9650 0.8475 2.0250 0.9075 ;
        RECT 1.8600 0.4650 1.9200 0.5250 ;
        RECT 1.7550 0.2250 1.8150 0.2850 ;
        RECT 1.7550 0.7200 1.8150 0.7800 ;
        RECT 1.6500 0.4650 1.7100 0.5250 ;
        RECT 1.5450 0.1275 1.6050 0.1875 ;
        RECT 1.5450 0.8250 1.6050 0.8850 ;
        RECT 1.4400 0.4800 1.5000 0.5400 ;
        RECT 1.3350 0.2250 1.3950 0.2850 ;
        RECT 1.3350 0.7575 1.3950 0.8175 ;
        RECT 1.2300 0.4800 1.2900 0.5400 ;
        RECT 1.1250 0.1200 1.1850 0.1800 ;
        RECT 1.1250 0.8700 1.1850 0.9300 ;
        RECT 1.0200 0.4875 1.0800 0.5475 ;
        RECT 0.8100 0.4200 0.8700 0.4800 ;
        RECT 0.8100 0.6600 0.8700 0.7200 ;
        RECT 0.7050 0.1725 0.7650 0.2325 ;
        RECT 0.7050 0.8325 0.7650 0.8925 ;
        RECT 0.5925 0.3450 0.6525 0.4050 ;
        RECT 0.3900 0.5700 0.4500 0.6300 ;
        RECT 0.3825 0.3300 0.4425 0.3900 ;
        RECT 0.2850 0.1350 0.3450 0.1950 ;
        RECT 0.2850 0.8625 0.3450 0.9225 ;
        RECT 0.1875 0.5400 0.2475 0.6000 ;
        RECT 0.0750 0.1575 0.1350 0.2175 ;
        RECT 0.0750 0.7950 0.1350 0.8550 ;
        LAYER M1 ;
        RECT 1.6575 0.4575 2.3700 0.5325 ;
        RECT 2.1525 0.1950 2.2575 0.3825 ;
        RECT 2.1675 0.6225 2.2425 0.8325 ;
        RECT 1.8225 0.6225 2.1675 0.7125 ;
        RECT 1.8375 0.2925 2.1525 0.3825 ;
        RECT 1.7325 0.1950 1.8375 0.3825 ;
        RECT 1.7475 0.6225 1.8225 0.8325 ;
        RECT 1.5825 0.2625 1.6575 0.7425 ;
        RECT 1.4175 0.2625 1.5825 0.3375 ;
        RECT 1.4100 0.6675 1.5825 0.7425 ;
        RECT 1.2600 0.4500 1.5000 0.5700 ;
        RECT 1.3350 0.1950 1.4175 0.3375 ;
        RECT 1.3350 0.6675 1.4100 0.8475 ;
        RECT 1.1850 0.2550 1.2600 0.7650 ;
        RECT 1.0200 0.2550 1.1850 0.3300 ;
        RECT 1.0425 0.6900 1.1850 0.7650 ;
        RECT 0.9675 0.4050 1.1100 0.6150 ;
        RECT 0.9675 0.6900 1.0425 0.9000 ;
        RECT 0.9450 0.1500 1.0200 0.3300 ;
        RECT 0.9450 0.4050 0.9675 0.5400 ;
        RECT 0.6750 0.8250 0.9675 0.9000 ;
        RECT 0.6825 0.1500 0.9450 0.2550 ;
        RECT 0.7875 0.6375 0.8925 0.7500 ;
        RECT 0.7875 0.3900 0.8700 0.5625 ;
        RECT 0.7200 0.4875 0.7875 0.5625 ;
        RECT 0.6000 0.6750 0.7875 0.7500 ;
        RECT 0.5700 0.4875 0.7200 0.6000 ;
        RECT 0.6075 0.3300 0.6825 0.4125 ;
        RECT 0.5175 0.1500 0.6075 0.4125 ;
        RECT 0.5400 0.6750 0.6000 0.7800 ;
        RECT 0.4800 0.5250 0.5700 0.6000 ;
        RECT 0.1425 0.7050 0.5400 0.7800 ;
        RECT 0.4875 0.1500 0.5175 0.2250 ;
        RECT 0.2925 0.5250 0.4800 0.6300 ;
        RECT 0.1650 0.3000 0.4425 0.4200 ;
        RECT 0.1875 0.5100 0.2925 0.6300 ;
        RECT 0.1125 0.1500 0.1650 0.4200 ;
        RECT 0.1125 0.7050 0.1425 0.9000 ;
        RECT 0.0375 0.1500 0.1125 0.9000 ;
    END
END MUX2N_0111


MACRO MUX2N_1000
    CLASS CORE ;
    FOREIGN MUX2N_1000 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.0900 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 5.4600 0.3150 5.6175 0.4350 ;
        RECT 5.4600 0.6150 5.6175 0.7350 ;
        RECT 5.1450 0.3150 5.4600 0.7350 ;
        RECT 4.9875 0.3150 5.1450 0.4350 ;
        RECT 4.9875 0.6150 5.1450 0.7350 ;
        VIA 5.4600 0.3750 VIA12_slot ;
        VIA 5.4600 0.6750 VIA12_slot ;
        VIA 5.1450 0.3750 VIA12_slot ;
        VIA 5.1450 0.6750 VIA12_slot ;
        END
    END ZN
    PIN S
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 2.8125 0.4125 3.5775 0.4875 ;
        RECT 2.7075 0.4125 2.8125 0.6075 ;
        VIA 3.4575 0.4500 VIA12_square ;
        VIA 2.7600 0.5175 VIA12_square ;
        END
    END S
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.5000 0.4575 1.6125 0.7875 ;
        RECT 0.9900 0.7125 1.5000 0.7875 ;
        VIA 1.5600 0.5400 VIA12_square ;
        END
    END I1
    PIN I0
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.6900 0.4350 0.8025 0.6375 ;
        RECT 0.1800 0.5625 0.6900 0.6375 ;
        VIA 0.7500 0.5175 VIA12_square ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 3.1200 -0.0750 6.0900 0.0750 ;
        RECT 2.9700 -0.0750 3.1200 0.2175 ;
        RECT 2.6850 -0.0750 2.9700 0.0750 ;
        RECT 2.5650 -0.0750 2.6850 0.2250 ;
        RECT 2.2650 -0.0750 2.5650 0.0750 ;
        RECT 2.1450 -0.0750 2.2650 0.2325 ;
        RECT 1.8450 -0.0750 2.1450 0.0750 ;
        RECT 1.7250 -0.0750 1.8450 0.2325 ;
        RECT 1.4250 -0.0750 1.7250 0.0750 ;
        RECT 1.3050 -0.0750 1.4250 0.2325 ;
        RECT 1.0050 -0.0750 1.3050 0.0750 ;
        RECT 0.8850 -0.0750 1.0050 0.2325 ;
        RECT 0.5775 -0.0750 0.8850 0.0750 ;
        RECT 0.4725 -0.0750 0.5775 0.2325 ;
        RECT 0.1650 -0.0750 0.4725 0.0750 ;
        RECT 0.0450 -0.0750 0.1650 0.2325 ;
        RECT 0.0000 -0.0750 0.0450 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 3.1050 0.9750 6.0900 1.1250 ;
        RECT 2.9850 0.8325 3.1050 1.1250 ;
        RECT 2.7000 0.9750 2.9850 1.1250 ;
        RECT 2.5500 0.8325 2.7000 1.1250 ;
        RECT 2.2650 0.9750 2.5500 1.1250 ;
        RECT 2.1450 0.8400 2.2650 1.1250 ;
        RECT 1.8450 0.9750 2.1450 1.1250 ;
        RECT 1.7250 0.8400 1.8450 1.1250 ;
        RECT 1.4250 0.9750 1.7250 1.1250 ;
        RECT 1.3050 0.8400 1.4250 1.1250 ;
        RECT 1.0050 0.9750 1.3050 1.1250 ;
        RECT 0.8850 0.8400 1.0050 1.1250 ;
        RECT 0.5850 0.9750 0.8850 1.1250 ;
        RECT 0.4650 0.8400 0.5850 1.1250 ;
        RECT 0.1650 0.9750 0.4650 1.1250 ;
        RECT 0.0450 0.8325 0.1650 1.1250 ;
        RECT 0.0000 0.9750 0.0450 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 5.9550 0.3075 6.0150 0.3675 ;
        RECT 5.9550 0.6750 6.0150 0.7350 ;
        RECT 5.8500 0.4950 5.9100 0.5550 ;
        RECT 5.7450 0.1575 5.8050 0.2175 ;
        RECT 5.7450 0.8325 5.8050 0.8925 ;
        RECT 5.6400 0.4950 5.7000 0.5550 ;
        RECT 5.5350 0.3225 5.5950 0.3825 ;
        RECT 5.5350 0.6750 5.5950 0.7350 ;
        RECT 5.4300 0.4950 5.4900 0.5550 ;
        RECT 5.3250 0.1575 5.3850 0.2175 ;
        RECT 5.3250 0.8325 5.3850 0.8925 ;
        RECT 5.2200 0.4950 5.2800 0.5550 ;
        RECT 5.1150 0.3225 5.1750 0.3825 ;
        RECT 5.1150 0.6750 5.1750 0.7350 ;
        RECT 5.0100 0.4950 5.0700 0.5550 ;
        RECT 4.9050 0.1575 4.9650 0.2175 ;
        RECT 4.9050 0.8325 4.9650 0.8925 ;
        RECT 4.8000 0.4950 4.8600 0.5550 ;
        RECT 4.6950 0.2625 4.7550 0.3225 ;
        RECT 4.6950 0.6750 4.7550 0.7350 ;
        RECT 4.5900 0.4800 4.6500 0.5400 ;
        RECT 4.4850 0.3000 4.5450 0.3600 ;
        RECT 4.4850 0.6675 4.5450 0.7275 ;
        RECT 4.3800 0.4800 4.4400 0.5400 ;
        RECT 4.2750 0.1575 4.3350 0.2175 ;
        RECT 4.2750 0.8325 4.3350 0.8925 ;
        RECT 4.1700 0.4800 4.2300 0.5400 ;
        RECT 4.0650 0.3000 4.1250 0.3600 ;
        RECT 4.0650 0.6675 4.1250 0.7275 ;
        RECT 3.9600 0.4800 4.0200 0.5400 ;
        RECT 3.8550 0.1575 3.9150 0.2175 ;
        RECT 3.8550 0.8325 3.9150 0.8925 ;
        RECT 3.7500 0.4800 3.8100 0.5400 ;
        RECT 3.6450 0.3000 3.7050 0.3600 ;
        RECT 3.6450 0.6825 3.7050 0.7425 ;
        RECT 3.5400 0.4800 3.6000 0.5400 ;
        RECT 3.4350 0.1875 3.4950 0.2475 ;
        RECT 3.4350 0.8025 3.4950 0.8625 ;
        RECT 3.2250 0.3075 3.2850 0.3675 ;
        RECT 3.2250 0.6900 3.2850 0.7500 ;
        RECT 3.1200 0.4875 3.1800 0.5475 ;
        RECT 3.0150 0.1575 3.0750 0.2175 ;
        RECT 3.0150 0.8325 3.0750 0.8925 ;
        RECT 2.9100 0.4875 2.9700 0.5475 ;
        RECT 2.8050 0.3075 2.8650 0.3675 ;
        RECT 2.8050 0.6900 2.8650 0.7500 ;
        RECT 2.7000 0.4875 2.7600 0.5475 ;
        RECT 2.5950 0.1425 2.6550 0.2025 ;
        RECT 2.5950 0.8325 2.6550 0.8925 ;
        RECT 2.4900 0.4875 2.5500 0.5475 ;
        RECT 2.3850 0.2925 2.4450 0.3525 ;
        RECT 2.3850 0.7200 2.4450 0.7800 ;
        RECT 2.2800 0.4875 2.3400 0.5475 ;
        RECT 2.1750 0.1650 2.2350 0.2250 ;
        RECT 2.1750 0.8475 2.2350 0.9075 ;
        RECT 2.0700 0.4875 2.1300 0.5475 ;
        RECT 1.9650 0.3075 2.0250 0.3675 ;
        RECT 1.9650 0.6900 2.0250 0.7500 ;
        RECT 1.8600 0.4875 1.9200 0.5475 ;
        RECT 1.7550 0.1650 1.8150 0.2250 ;
        RECT 1.7550 0.8475 1.8150 0.9075 ;
        RECT 1.6500 0.4875 1.7100 0.5475 ;
        RECT 1.5450 0.2925 1.6050 0.3525 ;
        RECT 1.5450 0.7350 1.6050 0.7950 ;
        RECT 1.4400 0.4875 1.5000 0.5475 ;
        RECT 1.3350 0.1650 1.3950 0.2250 ;
        RECT 1.3350 0.8475 1.3950 0.9075 ;
        RECT 1.2300 0.4875 1.2900 0.5475 ;
        RECT 1.1250 0.3075 1.1850 0.3675 ;
        RECT 1.1250 0.6900 1.1850 0.7500 ;
        RECT 1.0200 0.4875 1.0800 0.5475 ;
        RECT 0.9150 0.1650 0.9750 0.2250 ;
        RECT 0.9150 0.8475 0.9750 0.9075 ;
        RECT 0.8100 0.4875 0.8700 0.5475 ;
        RECT 0.7050 0.3075 0.7650 0.3675 ;
        RECT 0.7050 0.6900 0.7650 0.7500 ;
        RECT 0.6000 0.4875 0.6600 0.5475 ;
        RECT 0.4950 0.1500 0.5550 0.2100 ;
        RECT 0.4950 0.8475 0.5550 0.9075 ;
        RECT 0.3900 0.4875 0.4500 0.5475 ;
        RECT 0.2850 0.2925 0.3450 0.3525 ;
        RECT 0.2850 0.7350 0.3450 0.7950 ;
        RECT 0.1875 0.4875 0.2475 0.5475 ;
        RECT 0.0750 0.1650 0.1350 0.2250 ;
        RECT 0.0750 0.8325 0.1350 0.8925 ;
        LAYER M1 ;
        RECT 5.9250 0.2775 6.0450 0.4125 ;
        RECT 5.9400 0.6375 6.0225 0.7875 ;
        RECT 4.9200 0.4875 5.9700 0.5625 ;
        RECT 4.9875 0.6375 5.9400 0.7350 ;
        RECT 4.9875 0.3075 5.9250 0.4125 ;
        RECT 5.0325 0.1500 5.8575 0.2250 ;
        RECT 4.9875 0.8250 5.8350 0.9000 ;
        RECT 4.8675 0.1500 5.0325 0.2325 ;
        RECT 4.7625 0.3075 4.9875 0.3825 ;
        RECT 4.7175 0.6600 4.9875 0.7350 ;
        RECT 4.8225 0.8175 4.9875 0.9000 ;
        RECT 4.7250 0.4575 4.9200 0.5850 ;
        RECT 4.6875 0.1500 4.7625 0.3825 ;
        RECT 4.6425 0.6600 4.7175 0.9000 ;
        RECT 3.5100 0.1500 4.6875 0.2250 ;
        RECT 4.5450 0.4500 4.6500 0.5700 ;
        RECT 3.5025 0.8250 4.6425 0.9000 ;
        RECT 3.6150 0.3000 4.5750 0.3750 ;
        RECT 3.9825 0.6450 4.5675 0.7500 ;
        RECT 3.5100 0.4500 4.5450 0.5400 ;
        RECT 3.6150 0.6750 3.9825 0.7500 ;
        RECT 3.4050 0.1500 3.5100 0.2850 ;
        RECT 3.4050 0.3750 3.5100 0.5400 ;
        RECT 3.4275 0.7575 3.5025 0.9000 ;
        RECT 3.2550 0.3075 3.3300 0.7575 ;
        RECT 2.7675 0.3075 3.2550 0.3825 ;
        RECT 2.7675 0.6525 3.2550 0.7575 ;
        RECT 2.6625 0.4575 3.1800 0.5775 ;
        RECT 2.4225 0.4725 2.5800 0.5775 ;
        RECT 2.4525 0.3075 2.5575 0.3825 ;
        RECT 2.3775 0.2625 2.4525 0.3825 ;
        RECT 2.3775 0.6825 2.4525 0.8175 ;
        RECT 1.4400 0.4575 2.4225 0.5775 ;
        RECT 1.6125 0.3075 2.3775 0.3825 ;
        RECT 1.6125 0.6825 2.3775 0.7575 ;
        RECT 1.5375 0.2250 1.6125 0.3825 ;
        RECT 1.5375 0.6825 1.6125 0.8400 ;
        RECT 0.1875 0.4575 1.2900 0.5775 ;
        RECT 0.7725 0.3075 1.2675 0.3825 ;
        RECT 0.7725 0.6825 1.2675 0.7575 ;
        RECT 0.6975 0.2325 0.7725 0.3825 ;
        RECT 0.6975 0.6825 0.7725 0.8400 ;
        RECT 0.3525 0.3075 0.6975 0.3825 ;
        RECT 0.3525 0.6825 0.6975 0.7575 ;
        RECT 0.2775 0.2325 0.3525 0.3825 ;
        RECT 0.2775 0.6825 0.3525 0.8400 ;
        RECT 0.1125 0.3075 0.2775 0.3825 ;
        RECT 0.1125 0.6825 0.2775 0.7575 ;
        RECT 0.0375 0.3075 0.1125 0.7575 ;
        LAYER VIA1 ;
        RECT 4.9125 0.1575 4.9875 0.2325 ;
        RECT 4.8675 0.8175 4.9425 0.8925 ;
        RECT 4.7625 0.4800 4.8375 0.5550 ;
        RECT 4.0275 0.6675 4.1025 0.7425 ;
        RECT 3.8025 0.3000 3.8775 0.3750 ;
        RECT 3.2550 0.5625 3.3300 0.6375 ;
        RECT 2.4375 0.3075 2.5125 0.3825 ;
        RECT 2.0100 0.6825 2.0850 0.7575 ;
        RECT 1.9650 0.3075 2.0400 0.3825 ;
        RECT 1.1175 0.3075 1.1925 0.3825 ;
        LAYER M2 ;
        RECT 5.4900 0.3150 5.6175 0.4350 ;
        RECT 5.4900 0.6150 5.6175 0.7350 ;
        RECT 4.9875 0.3150 5.1150 0.4350 ;
        RECT 4.9875 0.6150 5.1150 0.7350 ;
        RECT 4.8675 0.1125 5.0325 0.2325 ;
        RECT 4.8225 0.8175 4.9875 0.9375 ;
        RECT 2.2950 0.1125 4.8675 0.1875 ;
        RECT 4.7625 0.4275 4.8375 0.6225 ;
        RECT 2.0850 0.8625 4.8225 0.9375 ;
        RECT 4.1175 0.4275 4.7625 0.5025 ;
        RECT 4.0125 0.6225 4.1250 0.7875 ;
        RECT 4.0425 0.4275 4.1175 0.5475 ;
        RECT 3.9375 0.4725 4.0425 0.5475 ;
        RECT 2.2950 0.7125 4.0125 0.7875 ;
        RECT 3.8625 0.4725 3.9375 0.6375 ;
        RECT 3.7575 0.2625 3.9225 0.3900 ;
        RECT 3.1950 0.5625 3.8625 0.6375 ;
        RECT 2.5275 0.2625 3.7575 0.3375 ;
        RECT 2.4225 0.2625 2.5275 0.4275 ;
        RECT 2.2200 0.1125 2.2950 0.7875 ;
        RECT 1.2075 0.1125 2.2200 0.1875 ;
        RECT 2.0100 0.3075 2.0850 0.9375 ;
        RECT 1.8975 0.3075 2.0100 0.3825 ;
        RECT 1.0950 0.1125 1.2075 0.4425 ;
    END
END MUX2N_1000


MACRO MUX2N_1010
    CLASS CORE ;
    FOREIGN MUX2N_1010 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.2600 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 0.9000 0.2625 1.1175 0.3375 ;
        RECT 0.9000 0.8625 0.9600 0.9375 ;
        RECT 0.8250 0.2625 0.9000 0.9375 ;
        RECT 0.4950 0.8625 0.8250 0.9375 ;
        VIA 1.0050 0.3000 VIA12_square ;
        VIA 0.8625 0.8325 VIA12_square ;
        END
    END ZN
    PIN S
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.1950 0.5625 0.6600 0.6375 ;
        VIA 0.3075 0.6000 VIA12_square ;
        END
    END S
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.1175 0.3675 1.2225 0.6825 ;
        RECT 1.0200 0.5625 1.1175 0.6825 ;
        END
    END I1
    PIN I0
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.1950 0.2625 0.6750 0.3375 ;
        VIA 0.5625 0.3000 VIA12_square ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.1925 -0.0750 1.2600 0.0750 ;
        RECT 1.1175 -0.0750 1.1925 0.2475 ;
        RECT 0.3750 -0.0750 1.1175 0.0750 ;
        RECT 0.2550 -0.0750 0.3750 0.2100 ;
        RECT 0.0000 -0.0750 0.2550 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.2000 0.9750 1.2600 1.1250 ;
        RECT 1.1250 0.8025 1.2000 1.1250 ;
        RECT 0.3750 0.9750 1.1250 1.1250 ;
        RECT 0.2550 0.8700 0.3750 1.1250 ;
        RECT 0.0000 0.9750 0.2550 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.1250 0.1575 1.1850 0.2175 ;
        RECT 1.1250 0.8325 1.1850 0.8925 ;
        RECT 1.0200 0.5925 1.0800 0.6525 ;
        RECT 0.8100 0.3600 0.8700 0.4200 ;
        RECT 0.8100 0.6450 0.8700 0.7050 ;
        RECT 0.7050 0.1725 0.7650 0.2325 ;
        RECT 0.7050 0.8175 0.7650 0.8775 ;
        RECT 0.5925 0.3450 0.6525 0.4050 ;
        RECT 0.3825 0.3150 0.4425 0.3750 ;
        RECT 0.3825 0.5550 0.4425 0.6150 ;
        RECT 0.2850 0.1350 0.3450 0.1950 ;
        RECT 0.2850 0.8700 0.3450 0.9300 ;
        RECT 0.1875 0.5550 0.2475 0.6150 ;
        RECT 0.0750 0.1575 0.1350 0.2175 ;
        RECT 0.0750 0.7950 0.1350 0.8550 ;
        LAYER M1 ;
        RECT 0.9675 0.1500 1.0425 0.3900 ;
        RECT 0.6675 0.7875 0.9900 0.9000 ;
        RECT 0.6825 0.1500 0.9675 0.2550 ;
        RECT 0.5925 0.6375 0.9000 0.7125 ;
        RECT 0.7875 0.3375 0.8925 0.5625 ;
        RECT 0.4425 0.4875 0.7875 0.5625 ;
        RECT 0.6075 0.3300 0.6825 0.4125 ;
        RECT 0.5175 0.1500 0.6075 0.4125 ;
        RECT 0.5175 0.6375 0.5925 0.7950 ;
        RECT 0.4875 0.1500 0.5175 0.2250 ;
        RECT 0.1425 0.7200 0.5175 0.7950 ;
        RECT 0.1650 0.2850 0.4425 0.4050 ;
        RECT 0.3525 0.4875 0.4425 0.6450 ;
        RECT 0.1875 0.5250 0.3525 0.6450 ;
        RECT 0.1125 0.1500 0.1650 0.4050 ;
        RECT 0.1125 0.7200 0.1425 0.9000 ;
        RECT 0.0375 0.1500 0.1125 0.9000 ;
    END
END MUX2N_1010


MACRO MUX2_0000
    CLASS CORE ;
    FOREIGN MUX2_0000 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.9900 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 3.4125 0.2775 3.5700 0.3975 ;
        RECT 3.4125 0.6525 3.5700 0.7725 ;
        RECT 3.0975 0.2775 3.4125 0.7725 ;
        RECT 2.9400 0.2775 3.0975 0.3975 ;
        RECT 2.9400 0.6525 3.0975 0.7725 ;
        VIA 3.4125 0.3375 VIA12_slot ;
        VIA 3.4125 0.7125 VIA12_slot ;
        VIA 3.0975 0.3375 VIA12_slot ;
        VIA 3.0975 0.7125 VIA12_slot ;
        END
    END Z
    PIN S
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.2825 0.5475 1.5825 0.6525 ;
        RECT 1.1175 0.4500 1.2825 0.6525 ;
        VIA 1.2000 0.4875 VIA12_square ;
        END
    END S
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.4425 0.4125 0.5475 0.6300 ;
        RECT 0.0675 0.4125 0.4425 0.4875 ;
        VIA 0.4950 0.5475 VIA12_square ;
        END
    END I1
    PIN I0
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.6375 0.4500 0.7425 0.7875 ;
        RECT 0.2175 0.7125 0.6375 0.7875 ;
        VIA 0.6900 0.5325 VIA12_square ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 3.9450 -0.0750 3.9900 0.0750 ;
        RECT 3.8250 -0.0750 3.9450 0.2925 ;
        RECT 3.5250 -0.0750 3.8250 0.0750 ;
        RECT 3.4050 -0.0750 3.5250 0.2025 ;
        RECT 3.1050 -0.0750 3.4050 0.0750 ;
        RECT 2.9850 -0.0750 3.1050 0.2025 ;
        RECT 2.6625 -0.0750 2.9850 0.0750 ;
        RECT 2.5875 -0.0750 2.6625 0.2475 ;
        RECT 1.0050 -0.0750 2.5875 0.0750 ;
        RECT 0.8850 -0.0750 1.0050 0.1875 ;
        RECT 0.5850 -0.0750 0.8850 0.0750 ;
        RECT 0.4650 -0.0750 0.5850 0.1875 ;
        RECT 0.1650 -0.0750 0.4650 0.0750 ;
        RECT 0.0450 -0.0750 0.1650 0.2175 ;
        RECT 0.0000 -0.0750 0.0450 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 3.9450 0.9750 3.9900 1.1250 ;
        RECT 3.8250 0.6600 3.9450 1.1250 ;
        RECT 3.5250 0.9750 3.8250 1.1250 ;
        RECT 3.4050 0.8475 3.5250 1.1250 ;
        RECT 3.1050 0.9750 3.4050 1.1250 ;
        RECT 2.9850 0.8475 3.1050 1.1250 ;
        RECT 2.6625 0.9750 2.9850 1.1250 ;
        RECT 2.5875 0.8025 2.6625 1.1250 ;
        RECT 0.9750 0.9750 2.5875 1.1250 ;
        RECT 0.8700 0.8400 0.9750 1.1250 ;
        RECT 0.5850 0.9750 0.8700 1.1250 ;
        RECT 0.4650 0.8625 0.5850 1.1250 ;
        RECT 0.1650 0.9750 0.4650 1.1250 ;
        RECT 0.0375 0.8325 0.1650 1.1250 ;
        RECT 0.0000 0.9750 0.0375 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 3.8550 0.2250 3.9150 0.2850 ;
        RECT 3.8550 0.6675 3.9150 0.7275 ;
        RECT 3.8550 0.8325 3.9150 0.8925 ;
        RECT 3.7500 0.4800 3.8100 0.5400 ;
        RECT 3.6450 0.3075 3.7050 0.3675 ;
        RECT 3.6450 0.6825 3.7050 0.7425 ;
        RECT 3.5400 0.4800 3.6000 0.5400 ;
        RECT 3.4350 0.1350 3.4950 0.1950 ;
        RECT 3.4350 0.8550 3.4950 0.9150 ;
        RECT 3.3300 0.4800 3.3900 0.5400 ;
        RECT 3.2250 0.3075 3.2850 0.3675 ;
        RECT 3.2250 0.6825 3.2850 0.7425 ;
        RECT 3.1200 0.4800 3.1800 0.5400 ;
        RECT 3.0150 0.1350 3.0750 0.1950 ;
        RECT 3.0150 0.8550 3.0750 0.9150 ;
        RECT 2.9100 0.4800 2.9700 0.5400 ;
        RECT 2.8050 0.3075 2.8650 0.3675 ;
        RECT 2.8050 0.6825 2.8650 0.7425 ;
        RECT 2.7000 0.4800 2.7600 0.5400 ;
        RECT 2.5950 0.1575 2.6550 0.2175 ;
        RECT 2.5950 0.8325 2.6550 0.8925 ;
        RECT 2.3850 0.1650 2.4450 0.2250 ;
        RECT 2.3850 0.8250 2.4450 0.8850 ;
        RECT 2.2725 0.4950 2.3325 0.5550 ;
        RECT 2.1750 0.3150 2.2350 0.3750 ;
        RECT 2.1750 0.6750 2.2350 0.7350 ;
        RECT 2.0775 0.4950 2.1375 0.5550 ;
        RECT 1.9650 0.1575 2.0250 0.2175 ;
        RECT 1.9650 0.8250 2.0250 0.8850 ;
        RECT 1.7550 0.1575 1.8150 0.2175 ;
        RECT 1.7550 0.8325 1.8150 0.8925 ;
        RECT 1.6500 0.4800 1.7100 0.5400 ;
        RECT 1.5450 0.3000 1.6050 0.3600 ;
        RECT 1.5450 0.6750 1.6050 0.7350 ;
        RECT 1.4325 0.4725 1.4925 0.5325 ;
        RECT 1.3350 0.1575 1.3950 0.2175 ;
        RECT 1.3350 0.8100 1.3950 0.8700 ;
        RECT 1.1250 0.2700 1.1850 0.3300 ;
        RECT 1.1250 0.8175 1.1850 0.8775 ;
        RECT 1.0275 0.4650 1.0875 0.5250 ;
        RECT 0.9150 0.1275 0.9750 0.1875 ;
        RECT 0.9150 0.8700 0.9750 0.9300 ;
        RECT 0.8025 0.4650 0.8625 0.5250 ;
        RECT 0.7050 0.2700 0.7650 0.3300 ;
        RECT 0.7050 0.7050 0.7650 0.7650 ;
        RECT 0.6075 0.4875 0.6675 0.5475 ;
        RECT 0.4950 0.1275 0.5550 0.1875 ;
        RECT 0.4950 0.8625 0.5550 0.9225 ;
        RECT 0.3900 0.4950 0.4500 0.5550 ;
        RECT 0.2850 0.2700 0.3450 0.3300 ;
        RECT 0.2850 0.7350 0.3450 0.7950 ;
        RECT 0.1875 0.4950 0.2475 0.5550 ;
        RECT 0.0750 0.1575 0.1350 0.2175 ;
        RECT 0.0750 0.8325 0.1350 0.8925 ;
        LAYER M1 ;
        RECT 2.4825 0.4725 3.8550 0.5475 ;
        RECT 2.7975 0.2775 3.7200 0.3975 ;
        RECT 2.7975 0.6525 3.7200 0.7725 ;
        RECT 2.4075 0.1500 2.4825 0.9000 ;
        RECT 1.3050 0.1500 2.4075 0.2250 ;
        RECT 1.4400 0.8250 2.4075 0.9000 ;
        RECT 2.2275 0.4650 2.3325 0.5925 ;
        RECT 2.1675 0.3075 2.3025 0.3825 ;
        RECT 1.9425 0.6675 2.3025 0.7425 ;
        RECT 2.0175 0.4875 2.2275 0.5925 ;
        RECT 1.9650 0.3075 2.1675 0.4125 ;
        RECT 1.8900 0.4875 1.9425 0.7425 ;
        RECT 1.8675 0.3000 1.8900 0.7425 ;
        RECT 1.8150 0.3000 1.8675 0.5625 ;
        RECT 1.4550 0.3000 1.8150 0.3750 ;
        RECT 1.5750 0.6450 1.7925 0.7500 ;
        RECT 1.6350 0.4500 1.7400 0.5700 ;
        RECT 1.4025 0.4500 1.6350 0.5325 ;
        RECT 1.5150 0.6150 1.5750 0.7500 ;
        RECT 1.3650 0.6150 1.5150 0.6900 ;
        RECT 1.3350 0.7800 1.4400 0.9000 ;
        RECT 0.9975 0.4500 1.4025 0.5250 ;
        RECT 1.3200 0.6000 1.3650 0.6900 ;
        RECT 0.9450 0.6000 1.3200 0.6750 ;
        RECT 1.0500 0.7500 1.2600 0.9000 ;
        RECT 1.0800 0.1650 1.1850 0.3750 ;
        RECT 0.9600 0.2700 1.0800 0.3750 ;
        RECT 0.8700 0.6000 0.9450 0.7650 ;
        RECT 0.7650 0.4425 0.8925 0.5250 ;
        RECT 0.8025 0.2625 0.8850 0.3675 ;
        RECT 0.6600 0.6900 0.8700 0.7650 ;
        RECT 0.6750 0.1500 0.8025 0.3675 ;
        RECT 0.6075 0.4425 0.7650 0.6150 ;
        RECT 0.3150 0.2625 0.5400 0.3375 ;
        RECT 0.4500 0.4650 0.5325 0.7125 ;
        RECT 0.1875 0.4650 0.4500 0.5850 ;
        RECT 0.2700 0.6825 0.3450 0.8325 ;
        RECT 0.2400 0.2625 0.3150 0.3900 ;
        RECT 0.1125 0.6825 0.2700 0.7575 ;
        RECT 0.1125 0.3150 0.2400 0.3900 ;
        RECT 0.0375 0.3150 0.1125 0.7575 ;
        LAYER VIA1 ;
        RECT 2.0625 0.5100 2.1375 0.5850 ;
        RECT 2.0100 0.3075 2.0850 0.3825 ;
        RECT 1.6725 0.6600 1.7475 0.7350 ;
        RECT 1.5000 0.3000 1.5750 0.3750 ;
        RECT 1.1250 0.7950 1.2000 0.8700 ;
        RECT 1.0200 0.2700 1.0950 0.3450 ;
        RECT 0.8175 0.6900 0.8925 0.7650 ;
        RECT 0.7350 0.2625 0.8100 0.3375 ;
        RECT 0.4200 0.2625 0.4950 0.3375 ;
        LAYER M2 ;
        RECT 3.4425 0.2775 3.5700 0.3975 ;
        RECT 3.4425 0.6525 3.5700 0.7725 ;
        RECT 2.9400 0.2775 3.0675 0.3975 ;
        RECT 2.9400 0.6525 3.0675 0.7725 ;
        RECT 2.0475 0.4650 2.1525 0.9375 ;
        RECT 1.8375 0.3075 2.1300 0.3825 ;
        RECT 1.2000 0.8625 2.0475 0.9375 ;
        RECT 1.7625 0.3075 1.8375 0.7800 ;
        RECT 1.6725 0.6150 1.7625 0.7800 ;
        RECT 1.5300 0.3000 1.6200 0.3750 ;
        RECT 1.4550 0.1125 1.5300 0.3750 ;
        RECT 0.5400 0.1125 1.4550 0.1875 ;
        RECT 1.1250 0.7425 1.2000 0.9375 ;
        RECT 1.0425 0.2700 1.1475 0.3450 ;
        RECT 1.0425 0.7425 1.1250 0.8175 ;
        RECT 0.9675 0.2700 1.0425 0.8175 ;
        RECT 0.8175 0.2625 0.8925 0.8100 ;
        RECT 0.6900 0.2625 0.8175 0.3375 ;
        RECT 0.4650 0.1125 0.5400 0.3375 ;
        RECT 0.3750 0.2625 0.4650 0.3375 ;
    END
END MUX2_0000


MACRO MUX2_0011
    CLASS CORE ;
    FOREIGN MUX2_0011 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.6800 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 1.5675 0.3075 1.6425 0.7425 ;
        RECT 1.4025 0.3075 1.5675 0.3825 ;
        RECT 1.4025 0.6675 1.5675 0.7425 ;
        RECT 1.3275 0.2175 1.4025 0.3825 ;
        RECT 1.3275 0.6675 1.4025 0.8325 ;
        END
    END Z
    PIN S
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.5025 0.7125 0.9225 0.7875 ;
        RECT 0.3975 0.4875 0.5025 0.7875 ;
        VIA 0.4500 0.5625 VIA12_square ;
        END
    END S
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.6525 0.4125 1.1175 0.4875 ;
        VIA 1.0200 0.4500 VIA12_square ;
        END
    END I1
    PIN I0
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.4275 0.2625 0.8925 0.3375 ;
        VIA 0.5625 0.3000 VIA12_square ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.6350 -0.0750 1.6800 0.0750 ;
        RECT 1.5150 -0.0750 1.6350 0.2250 ;
        RECT 1.2150 -0.0750 1.5150 0.0750 ;
        RECT 1.0950 -0.0750 1.2150 0.1800 ;
        RECT 0.3750 -0.0750 1.0950 0.0750 ;
        RECT 0.2550 -0.0750 0.3750 0.1800 ;
        RECT 0.0000 -0.0750 0.2550 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.6350 0.9750 1.6800 1.1250 ;
        RECT 1.5150 0.8250 1.6350 1.1250 ;
        RECT 1.2300 0.9750 1.5150 1.1250 ;
        RECT 1.1250 0.8400 1.2300 1.1250 ;
        RECT 0.3750 0.9750 1.1250 1.1250 ;
        RECT 0.2550 0.8625 0.3750 1.1250 ;
        RECT 0.0000 0.9750 0.2550 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.5450 0.1575 1.6050 0.2175 ;
        RECT 1.5450 0.8325 1.6050 0.8925 ;
        RECT 1.4325 0.4875 1.4925 0.5475 ;
        RECT 1.3350 0.2700 1.3950 0.3300 ;
        RECT 1.3350 0.7200 1.3950 0.7800 ;
        RECT 1.2300 0.4875 1.2900 0.5475 ;
        RECT 1.1250 0.1200 1.1850 0.1800 ;
        RECT 1.1250 0.8700 1.1850 0.9300 ;
        RECT 1.0200 0.4875 1.0800 0.5475 ;
        RECT 0.8100 0.6600 0.8700 0.7200 ;
        RECT 0.8025 0.4200 0.8625 0.4800 ;
        RECT 0.7050 0.1725 0.7650 0.2325 ;
        RECT 0.7050 0.8325 0.7650 0.8925 ;
        RECT 0.5925 0.3450 0.6525 0.4050 ;
        RECT 0.3825 0.3150 0.4425 0.3750 ;
        RECT 0.3825 0.5550 0.4425 0.6150 ;
        RECT 0.2850 0.1200 0.3450 0.1800 ;
        RECT 0.2850 0.8700 0.3450 0.9300 ;
        RECT 0.1875 0.5250 0.2475 0.5850 ;
        RECT 0.0750 0.7950 0.1350 0.8550 ;
        RECT 0.0750 0.1575 0.1350 0.2175 ;
        LAYER M1 ;
        RECT 1.2525 0.4575 1.4925 0.5775 ;
        RECT 1.1775 0.2550 1.2525 0.7650 ;
        RECT 1.0200 0.2550 1.1775 0.3300 ;
        RECT 1.0500 0.6900 1.1775 0.7650 ;
        RECT 0.9675 0.4050 1.1025 0.6150 ;
        RECT 0.9750 0.6900 1.0500 0.9000 ;
        RECT 0.9450 0.1500 1.0200 0.3300 ;
        RECT 0.6750 0.8250 0.9750 0.9000 ;
        RECT 0.9375 0.4050 0.9675 0.5400 ;
        RECT 0.6825 0.1500 0.9450 0.2550 ;
        RECT 0.7875 0.6375 0.8925 0.7500 ;
        RECT 0.7875 0.3900 0.8625 0.5625 ;
        RECT 0.7200 0.4875 0.7875 0.5625 ;
        RECT 0.6150 0.6750 0.7875 0.7500 ;
        RECT 0.6525 0.4875 0.7200 0.6000 ;
        RECT 0.6075 0.3300 0.6825 0.4125 ;
        RECT 0.4725 0.5250 0.6525 0.6000 ;
        RECT 0.5475 0.6750 0.6150 0.7650 ;
        RECT 0.5925 0.1500 0.6075 0.4125 ;
        RECT 0.5175 0.1500 0.5925 0.4200 ;
        RECT 0.1425 0.6900 0.5475 0.7650 ;
        RECT 0.5025 0.1500 0.5175 0.2250 ;
        RECT 0.2925 0.5250 0.4725 0.6150 ;
        RECT 0.3375 0.2850 0.4425 0.4050 ;
        RECT 0.1650 0.3300 0.3375 0.4050 ;
        RECT 0.1875 0.4800 0.2925 0.6150 ;
        RECT 0.1125 0.1500 0.1650 0.4050 ;
        RECT 0.1125 0.6900 0.1425 0.9000 ;
        RECT 0.0375 0.1500 0.1125 0.9000 ;
    END
END MUX2_0011


MACRO MUX2_0111
    CLASS CORE ;
    FOREIGN MUX2_0111 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.1500 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 2.4675 0.2625 2.7825 0.7725 ;
        VIA 2.6250 0.3225 VIA12_slot ;
        VIA 2.6250 0.7125 VIA12_slot ;
        END
    END Z
    PIN S
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.2450 0.3525 1.4175 0.4575 ;
        RECT 1.1700 0.1125 1.2450 0.4575 ;
        RECT 0.4275 0.1125 1.1700 0.1875 ;
        RECT 0.4275 0.5250 0.5475 0.6000 ;
        RECT 0.3525 0.1125 0.4275 0.6000 ;
        VIA 1.3425 0.4050 VIA12_square ;
        VIA 0.4350 0.5625 VIA12_square ;
        END
    END S
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 2.0850 0.8625 2.4000 0.9375 ;
        RECT 2.0100 0.4125 2.0850 0.9375 ;
        RECT 1.6950 0.4125 2.0100 0.4875 ;
        VIA 2.0475 0.5025 VIA12_square ;
        END
    END I1
    PIN I0
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.0125 0.2625 1.0875 0.6075 ;
        RECT 0.5475 0.2625 1.0125 0.3375 ;
        VIA 1.0500 0.5250 VIA12_square ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 3.0825 -0.0750 3.1500 0.0750 ;
        RECT 3.0075 -0.0750 3.0825 0.2625 ;
        RECT 2.6850 -0.0750 3.0075 0.0750 ;
        RECT 2.5650 -0.0750 2.6850 0.1950 ;
        RECT 2.2425 -0.0750 2.5650 0.0750 ;
        RECT 2.1675 -0.0750 2.2425 0.2475 ;
        RECT 1.8450 -0.0750 2.1675 0.0750 ;
        RECT 1.7250 -0.0750 1.8450 0.2250 ;
        RECT 0.7950 -0.0750 1.7250 0.0750 ;
        RECT 0.6750 -0.0750 0.7950 0.2175 ;
        RECT 0.3750 -0.0750 0.6750 0.0750 ;
        RECT 0.2550 -0.0750 0.3750 0.2250 ;
        RECT 0.0000 -0.0750 0.2550 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 3.0975 0.9750 3.1500 1.1250 ;
        RECT 2.9925 0.6375 3.0975 1.1250 ;
        RECT 2.6850 0.9750 2.9925 1.1250 ;
        RECT 2.5650 0.8400 2.6850 1.1250 ;
        RECT 2.2650 0.9750 2.5650 1.1250 ;
        RECT 2.1450 0.6600 2.2650 1.1250 ;
        RECT 1.8375 0.9750 2.1450 1.1250 ;
        RECT 1.7325 0.7800 1.8375 1.1250 ;
        RECT 0.7950 0.9750 1.7325 1.1250 ;
        RECT 0.6750 0.8325 0.7950 1.1250 ;
        RECT 0.3600 0.9750 0.6750 1.1250 ;
        RECT 0.2850 0.7950 0.3600 1.1250 ;
        RECT 0.0000 0.9750 0.2850 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 3.0150 0.1725 3.0750 0.2325 ;
        RECT 3.0150 0.6675 3.0750 0.7275 ;
        RECT 3.0150 0.8325 3.0750 0.8925 ;
        RECT 2.9100 0.4800 2.9700 0.5400 ;
        RECT 2.8050 0.2925 2.8650 0.3525 ;
        RECT 2.8050 0.6825 2.8650 0.7425 ;
        RECT 2.7000 0.4800 2.7600 0.5400 ;
        RECT 2.5950 0.1275 2.6550 0.1875 ;
        RECT 2.5950 0.8550 2.6550 0.9150 ;
        RECT 2.4900 0.4800 2.5500 0.5400 ;
        RECT 2.3850 0.2925 2.4450 0.3525 ;
        RECT 2.3850 0.6825 2.4450 0.7425 ;
        RECT 2.2800 0.4800 2.3400 0.5400 ;
        RECT 2.1750 0.1575 2.2350 0.2175 ;
        RECT 2.1750 0.6675 2.2350 0.7275 ;
        RECT 2.1750 0.8325 2.2350 0.8925 ;
        RECT 2.0625 0.4725 2.1225 0.5325 ;
        RECT 1.9650 0.2850 2.0250 0.3450 ;
        RECT 1.9650 0.6675 2.0250 0.7275 ;
        RECT 1.8600 0.4725 1.9200 0.5325 ;
        RECT 1.7550 0.1575 1.8150 0.2175 ;
        RECT 1.7550 0.8025 1.8150 0.8625 ;
        RECT 1.5450 0.1800 1.6050 0.2400 ;
        RECT 1.5450 0.8100 1.6050 0.8700 ;
        RECT 1.4400 0.3600 1.5000 0.4200 ;
        RECT 1.4400 0.6000 1.5000 0.6600 ;
        RECT 1.3350 0.1650 1.3950 0.2250 ;
        RECT 1.3350 0.8175 1.3950 0.8775 ;
        RECT 1.1250 0.1725 1.1850 0.2325 ;
        RECT 1.1250 0.8175 1.1850 0.8775 ;
        RECT 1.0200 0.4950 1.0800 0.5550 ;
        RECT 0.9150 0.2025 0.9750 0.2625 ;
        RECT 0.9150 0.6900 0.9750 0.7500 ;
        RECT 0.8100 0.5100 0.8700 0.5700 ;
        RECT 0.7050 0.1575 0.7650 0.2175 ;
        RECT 0.7050 0.8325 0.7650 0.8925 ;
        RECT 0.6000 0.5100 0.6600 0.5700 ;
        RECT 0.4950 0.1725 0.5550 0.2325 ;
        RECT 0.4950 0.7875 0.5550 0.8475 ;
        RECT 0.3900 0.3600 0.4500 0.4200 ;
        RECT 0.3900 0.6000 0.4500 0.6600 ;
        RECT 0.2850 0.1575 0.3450 0.2175 ;
        RECT 0.2850 0.8250 0.3450 0.8850 ;
        RECT 0.1875 0.5550 0.2475 0.6150 ;
        RECT 0.0750 0.2025 0.1350 0.2625 ;
        RECT 0.0750 0.7725 0.1350 0.8325 ;
        LAYER M1 ;
        RECT 2.2200 0.4575 3.0075 0.5625 ;
        RECT 2.3550 0.2700 2.8950 0.3750 ;
        RECT 2.3550 0.6600 2.8875 0.7650 ;
        RECT 1.8375 0.4500 2.1450 0.5550 ;
        RECT 1.9575 0.2550 2.0325 0.3750 ;
        RECT 1.9575 0.6300 2.0325 0.7575 ;
        RECT 1.6500 0.3000 1.9575 0.3750 ;
        RECT 1.6575 0.6300 1.9575 0.7050 ;
        RECT 1.5825 0.6300 1.6575 0.9000 ;
        RECT 1.5750 0.1500 1.6500 0.3750 ;
        RECT 1.5450 0.7800 1.5825 0.9000 ;
        RECT 1.5450 0.1500 1.5750 0.2700 ;
        RECT 1.2900 0.5550 1.5075 0.7050 ;
        RECT 1.2900 0.3300 1.5000 0.4800 ;
        RECT 1.1025 0.1500 1.4700 0.2550 ;
        RECT 1.1025 0.7950 1.4700 0.9000 ;
        RECT 1.0125 0.4425 1.2150 0.6075 ;
        RECT 0.6000 0.6825 1.0050 0.7575 ;
        RECT 0.9075 0.1725 0.9825 0.3675 ;
        RECT 0.7425 0.4425 0.9375 0.6075 ;
        RECT 0.6000 0.2925 0.9075 0.3675 ;
        RECT 0.5925 0.4800 0.6675 0.6000 ;
        RECT 0.5250 0.1500 0.6000 0.3675 ;
        RECT 0.5250 0.6825 0.6000 0.8775 ;
        RECT 0.4500 0.5250 0.5925 0.6000 ;
        RECT 0.4725 0.1500 0.5250 0.2550 ;
        RECT 0.4875 0.7575 0.5250 0.8775 ;
        RECT 0.3150 0.3300 0.4500 0.4500 ;
        RECT 0.3450 0.5250 0.4500 0.6900 ;
        RECT 0.1875 0.5250 0.3450 0.6450 ;
        RECT 0.1575 0.3300 0.3150 0.4050 ;
        RECT 0.1125 0.7275 0.2100 0.8925 ;
        RECT 0.1125 0.1800 0.1575 0.4050 ;
        RECT 0.0375 0.1800 0.1125 0.8925 ;
        LAYER VIA1 ;
        RECT 2.2575 0.4725 2.3325 0.5475 ;
        RECT 1.3575 0.1650 1.4325 0.2400 ;
        RECT 1.3575 0.8100 1.4325 0.8850 ;
        RECT 1.3050 0.5925 1.3800 0.6675 ;
        RECT 0.7875 0.4875 0.8625 0.5625 ;
        RECT 0.1350 0.7725 0.2100 0.8475 ;
        LAYER M2 ;
        RECT 2.3025 0.4275 2.3475 0.5925 ;
        RECT 2.2275 0.2625 2.3025 0.5925 ;
        RECT 1.5750 0.2625 2.2275 0.3375 ;
        RECT 1.5000 0.1500 1.5750 0.8700 ;
        RECT 1.3200 0.1500 1.5000 0.2550 ;
        RECT 1.4700 0.7950 1.5000 0.8700 ;
        RECT 1.3200 0.7950 1.4700 0.9000 ;
        RECT 1.2450 0.5775 1.4175 0.6825 ;
        RECT 1.1700 0.5775 1.2450 0.8475 ;
        RECT 0.8775 0.7725 1.1700 0.8475 ;
        RECT 0.7725 0.4425 0.8775 0.8475 ;
        RECT 0.0600 0.7725 0.7725 0.8475 ;
    END
END MUX2_0111


MACRO MUX2_1000
    CLASS CORE ;
    FOREIGN MUX2_1000 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.4700 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 1.3575 0.1500 1.4325 0.9000 ;
        RECT 1.3275 0.1500 1.3575 0.3825 ;
        RECT 1.3275 0.6675 1.3575 0.9000 ;
        END
    END Z
    PIN S
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.5025 0.7125 0.9225 0.7875 ;
        RECT 0.3975 0.4875 0.5025 0.7875 ;
        VIA 0.4500 0.5625 VIA12_square ;
        END
    END S
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.6525 0.4125 1.1175 0.4875 ;
        VIA 1.0200 0.4500 VIA12_square ;
        END
    END I1
    PIN I0
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.4275 0.2625 0.8925 0.3375 ;
        VIA 0.5625 0.3000 VIA12_square ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.2150 -0.0750 1.4700 0.0750 ;
        RECT 1.0950 -0.0750 1.2150 0.1800 ;
        RECT 0.3750 -0.0750 1.0950 0.0750 ;
        RECT 0.2550 -0.0750 0.3750 0.2100 ;
        RECT 0.0000 -0.0750 0.2550 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.2300 0.9750 1.4700 1.1250 ;
        RECT 1.1250 0.8400 1.2300 1.1250 ;
        RECT 0.3750 0.9750 1.1250 1.1250 ;
        RECT 0.2550 0.8400 0.3750 1.1250 ;
        RECT 0.0000 0.9750 0.2550 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.3350 0.1800 1.3950 0.2400 ;
        RECT 1.3350 0.8100 1.3950 0.8700 ;
        RECT 1.2225 0.4800 1.2825 0.5400 ;
        RECT 1.1250 0.1200 1.1850 0.1800 ;
        RECT 1.1250 0.8700 1.1850 0.9300 ;
        RECT 1.0200 0.4875 1.0800 0.5475 ;
        RECT 0.8100 0.6600 0.8700 0.7200 ;
        RECT 0.8025 0.4200 0.8625 0.4800 ;
        RECT 0.7050 0.1725 0.7650 0.2325 ;
        RECT 0.7050 0.8325 0.7650 0.8925 ;
        RECT 0.5925 0.3450 0.6525 0.4050 ;
        RECT 0.3825 0.3150 0.4425 0.3750 ;
        RECT 0.3825 0.5550 0.4425 0.6150 ;
        RECT 0.1875 0.5250 0.2475 0.5850 ;
        RECT 0.0750 0.1575 0.1350 0.2175 ;
        RECT 0.0750 0.8175 0.1350 0.8775 ;
        RECT 0.2850 0.1350 0.3450 0.1950 ;
        RECT 0.2850 0.8475 0.3450 0.9075 ;
        LAYER M1 ;
        RECT 1.2525 0.4500 1.2825 0.5700 ;
        RECT 1.1775 0.2550 1.2525 0.7650 ;
        RECT 1.0200 0.2550 1.1775 0.3300 ;
        RECT 1.0500 0.6900 1.1775 0.7650 ;
        RECT 0.9675 0.4050 1.1025 0.6150 ;
        RECT 0.9750 0.6900 1.0500 0.9000 ;
        RECT 0.9450 0.1500 1.0200 0.3300 ;
        RECT 0.6750 0.8250 0.9750 0.9000 ;
        RECT 0.9375 0.4050 0.9675 0.5400 ;
        RECT 0.6825 0.1500 0.9450 0.2550 ;
        RECT 0.7875 0.6375 0.8925 0.7500 ;
        RECT 0.7875 0.3900 0.8625 0.5625 ;
        RECT 0.7200 0.4875 0.7875 0.5625 ;
        RECT 0.6150 0.6750 0.7875 0.7500 ;
        RECT 0.6525 0.4875 0.7200 0.6000 ;
        RECT 0.6075 0.3300 0.6825 0.4125 ;
        RECT 0.4725 0.5250 0.6525 0.6000 ;
        RECT 0.5475 0.6750 0.6150 0.7650 ;
        RECT 0.5925 0.1500 0.6075 0.4125 ;
        RECT 0.5175 0.1500 0.5925 0.4200 ;
        RECT 0.1575 0.6900 0.5475 0.7650 ;
        RECT 0.5025 0.1500 0.5175 0.2250 ;
        RECT 0.2925 0.5250 0.4725 0.6150 ;
        RECT 0.3375 0.2850 0.4425 0.4050 ;
        RECT 0.1650 0.3300 0.3375 0.4050 ;
        RECT 0.1875 0.4800 0.2925 0.6150 ;
        RECT 0.1125 0.1500 0.1650 0.4050 ;
        RECT 0.1125 0.6900 0.1575 0.9000 ;
        RECT 0.0375 0.1500 0.1125 0.9000 ;
    END
END MUX2_1000


MACRO MUX2_1010
    CLASS CORE ;
    FOREIGN MUX2_1010 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.4700 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 1.3575 0.2025 1.4325 0.8325 ;
        RECT 1.3275 0.2025 1.3575 0.3825 ;
        RECT 1.3275 0.6675 1.3575 0.8325 ;
        END
    END Z
    PIN S
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.5025 0.7125 0.9225 0.7875 ;
        RECT 0.3975 0.4875 0.5025 0.7875 ;
        VIA 0.4500 0.5625 VIA12_square ;
        END
    END S
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.6525 0.4125 1.1175 0.4875 ;
        VIA 1.0200 0.4500 VIA12_square ;
        END
    END I1
    PIN I0
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.4275 0.2625 0.8925 0.3375 ;
        VIA 0.5625 0.3000 VIA12_square ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.2150 -0.0750 1.4700 0.0750 ;
        RECT 1.0950 -0.0750 1.2150 0.1800 ;
        RECT 0.3750 -0.0750 1.0950 0.0750 ;
        RECT 0.2550 -0.0750 0.3750 0.2025 ;
        RECT 0.0000 -0.0750 0.2550 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.2300 0.9750 1.4700 1.1250 ;
        RECT 1.1250 0.8400 1.2300 1.1250 ;
        RECT 0.3750 0.9750 1.1250 1.1250 ;
        RECT 0.2550 0.8400 0.3750 1.1250 ;
        RECT 0.0000 0.9750 0.2550 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.3350 0.2775 1.3950 0.3375 ;
        RECT 1.3350 0.7200 1.3950 0.7800 ;
        RECT 1.2225 0.4800 1.2825 0.5400 ;
        RECT 1.1250 0.1200 1.1850 0.1800 ;
        RECT 1.1250 0.8700 1.1850 0.9300 ;
        RECT 1.0200 0.4875 1.0800 0.5475 ;
        RECT 0.8100 0.6600 0.8700 0.7200 ;
        RECT 0.8025 0.4200 0.8625 0.4800 ;
        RECT 0.7050 0.1725 0.7650 0.2325 ;
        RECT 0.7050 0.8325 0.7650 0.8925 ;
        RECT 0.5925 0.3450 0.6525 0.4050 ;
        RECT 0.3825 0.3150 0.4425 0.3750 ;
        RECT 0.3825 0.5550 0.4425 0.6150 ;
        RECT 0.1875 0.5250 0.2475 0.5850 ;
        RECT 0.0750 0.1575 0.1350 0.2175 ;
        RECT 0.0750 0.7950 0.1350 0.8550 ;
        RECT 0.2850 0.1350 0.3450 0.1950 ;
        RECT 0.2850 0.8550 0.3450 0.9150 ;
        LAYER M1 ;
        RECT 1.2525 0.4500 1.2825 0.5700 ;
        RECT 1.1775 0.2550 1.2525 0.7650 ;
        RECT 1.0200 0.2550 1.1775 0.3300 ;
        RECT 1.0500 0.6900 1.1775 0.7650 ;
        RECT 0.9675 0.4050 1.1025 0.6150 ;
        RECT 0.9750 0.6900 1.0500 0.9000 ;
        RECT 0.9450 0.1500 1.0200 0.3300 ;
        RECT 0.6750 0.8250 0.9750 0.9000 ;
        RECT 0.9375 0.4050 0.9675 0.5400 ;
        RECT 0.6825 0.1500 0.9450 0.2550 ;
        RECT 0.7875 0.6375 0.8925 0.7500 ;
        RECT 0.7875 0.3900 0.8625 0.5625 ;
        RECT 0.7200 0.4875 0.7875 0.5625 ;
        RECT 0.6150 0.6750 0.7875 0.7500 ;
        RECT 0.6525 0.4875 0.7200 0.6000 ;
        RECT 0.6075 0.3300 0.6825 0.4125 ;
        RECT 0.4725 0.5250 0.6525 0.6000 ;
        RECT 0.5475 0.6750 0.6150 0.7650 ;
        RECT 0.5925 0.1500 0.6075 0.4125 ;
        RECT 0.5175 0.1500 0.5925 0.4200 ;
        RECT 0.1425 0.6900 0.5475 0.7650 ;
        RECT 0.5025 0.1500 0.5175 0.2250 ;
        RECT 0.2925 0.5250 0.4725 0.6150 ;
        RECT 0.3375 0.2850 0.4425 0.4050 ;
        RECT 0.1650 0.3300 0.3375 0.4050 ;
        RECT 0.1875 0.4800 0.2925 0.6150 ;
        RECT 0.1125 0.1500 0.1650 0.4050 ;
        RECT 0.1125 0.6900 0.1425 0.9000 ;
        RECT 0.0375 0.1500 0.1125 0.9000 ;
    END
END MUX2_1010


MACRO MUX3N_0011
    CLASS CORE ;
    FOREIGN MUX3N_0011 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.3600 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 3.2475 0.3000 3.3225 0.7425 ;
        RECT 3.0825 0.3000 3.2475 0.3825 ;
        RECT 3.0825 0.6675 3.2475 0.7425 ;
        RECT 3.0075 0.2175 3.0825 0.3825 ;
        RECT 3.0075 0.6675 3.0825 0.8325 ;
        END
    END ZN
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.9125 0.1125 2.3775 0.1875 ;
        RECT 1.8375 0.1125 1.9125 0.6000 ;
        VIA 1.8750 0.5175 VIA12_square ;
        END
    END S1
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.4275 0.1125 0.7200 0.1875 ;
        RECT 0.4275 0.2625 0.6450 0.3375 ;
        RECT 0.3525 0.1125 0.4275 0.6900 ;
        RECT 0.1800 0.1125 0.3525 0.1875 ;
        VIA 0.5625 0.3000 VIA12_square ;
        VIA 0.3900 0.6075 VIA12_square ;
        END
    END S0
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 2.1975 0.5625 2.6625 0.6375 ;
        VIA 2.3250 0.6000 VIA12_square ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.9525 0.5625 1.4175 0.6375 ;
        VIA 1.0725 0.6000 VIA12_square ;
        END
    END I1
    PIN I0
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.6375 0.4125 1.1175 0.4875 ;
        RECT 0.5325 0.4125 0.6375 0.7500 ;
        VIA 0.5850 0.6675 VIA12_square ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 3.3150 -0.0750 3.3600 0.0750 ;
        RECT 3.1950 -0.0750 3.3150 0.2250 ;
        RECT 2.8725 -0.0750 3.1950 0.0750 ;
        RECT 2.7975 -0.0750 2.8725 0.3000 ;
        RECT 2.4750 -0.0750 2.7975 0.0750 ;
        RECT 2.3550 -0.0750 2.4750 0.1800 ;
        RECT 1.1850 -0.0750 2.3550 0.0750 ;
        RECT 1.0800 -0.0750 1.1850 0.2475 ;
        RECT 0.3750 -0.0750 1.0800 0.0750 ;
        RECT 0.2550 -0.0750 0.3750 0.1800 ;
        RECT 0.0000 -0.0750 0.2550 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 3.3150 0.9750 3.3600 1.1250 ;
        RECT 3.1950 0.8250 3.3150 1.1250 ;
        RECT 2.8875 0.9750 3.1950 1.1250 ;
        RECT 2.7825 0.6450 2.8875 1.1250 ;
        RECT 2.4750 0.9750 2.7825 1.1250 ;
        RECT 2.3550 0.7875 2.4750 1.1250 ;
        RECT 1.2000 0.9750 2.3550 1.1250 ;
        RECT 1.1250 0.7875 1.2000 1.1250 ;
        RECT 0.3750 0.9750 1.1250 1.1250 ;
        RECT 0.2550 0.7650 0.3750 1.1250 ;
        RECT 0.0000 0.9750 0.2550 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 3.2250 0.1575 3.2850 0.2175 ;
        RECT 3.2250 0.8325 3.2850 0.8925 ;
        RECT 3.1125 0.4875 3.1725 0.5475 ;
        RECT 3.0150 0.2700 3.0750 0.3300 ;
        RECT 3.0150 0.7200 3.0750 0.7800 ;
        RECT 2.9100 0.4800 2.9700 0.5400 ;
        RECT 2.8050 0.2100 2.8650 0.2700 ;
        RECT 2.8050 0.6675 2.8650 0.7275 ;
        RECT 2.8050 0.8325 2.8650 0.8925 ;
        RECT 2.5950 0.2700 2.6550 0.3300 ;
        RECT 2.5950 0.7500 2.6550 0.8100 ;
        RECT 2.4825 0.4800 2.5425 0.5400 ;
        RECT 2.3850 0.1200 2.4450 0.1800 ;
        RECT 2.3850 0.8175 2.4450 0.8775 ;
        RECT 2.2800 0.4500 2.3400 0.5100 ;
        RECT 2.0700 0.3975 2.1300 0.4575 ;
        RECT 2.0700 0.6375 2.1300 0.6975 ;
        RECT 1.9650 0.1650 2.0250 0.2250 ;
        RECT 1.9650 0.8100 2.0250 0.8700 ;
        RECT 1.8600 0.4875 1.9200 0.5475 ;
        RECT 1.7550 0.1650 1.8150 0.2250 ;
        RECT 1.7550 0.8175 1.8150 0.8775 ;
        RECT 1.6500 0.3375 1.7100 0.3975 ;
        RECT 1.5450 0.1650 1.6050 0.2250 ;
        RECT 1.3350 0.3075 1.3950 0.3675 ;
        RECT 1.3350 0.7350 1.3950 0.7950 ;
        RECT 1.2300 0.4875 1.2900 0.5475 ;
        RECT 1.1250 0.1575 1.1850 0.2175 ;
        RECT 1.1250 0.8175 1.1850 0.8775 ;
        RECT 1.0200 0.4650 1.0800 0.5250 ;
        RECT 0.8100 0.3600 0.8700 0.4200 ;
        RECT 0.8100 0.6000 0.8700 0.6600 ;
        RECT 0.7050 0.1725 0.7650 0.2325 ;
        RECT 0.7050 0.8325 0.7650 0.8925 ;
        RECT 0.6000 0.5700 0.6600 0.6300 ;
        RECT 0.3900 0.3600 0.4500 0.4200 ;
        RECT 0.3900 0.6000 0.4500 0.6600 ;
        RECT 0.2850 0.1200 0.3450 0.1800 ;
        RECT 0.2850 0.7950 0.3450 0.8550 ;
        RECT 0.1875 0.5025 0.2475 0.5625 ;
        RECT 0.0750 0.1950 0.1350 0.2550 ;
        RECT 0.0750 0.7725 0.1350 0.8325 ;
        LAYER M1 ;
        RECT 3.0675 0.4575 3.1725 0.5775 ;
        RECT 2.6925 0.4575 3.0675 0.5475 ;
        RECT 2.6175 0.2175 2.6925 0.8400 ;
        RECT 2.5875 0.2175 2.6175 0.3825 ;
        RECT 2.5875 0.7200 2.6175 0.8400 ;
        RECT 2.5125 0.4500 2.5425 0.5700 ;
        RECT 2.4375 0.2625 2.5125 0.5700 ;
        RECT 2.2800 0.2625 2.4375 0.3375 ;
        RECT 2.2725 0.4125 2.3625 0.6825 ;
        RECT 2.2050 0.1500 2.2800 0.3375 ;
        RECT 2.2050 0.4125 2.2725 0.5625 ;
        RECT 1.9125 0.7800 2.2275 0.9000 ;
        RECT 1.8825 0.1500 2.2050 0.2400 ;
        RECT 1.4025 0.6300 2.1675 0.7050 ;
        RECT 2.0250 0.3675 2.1300 0.5550 ;
        RECT 1.2675 0.4800 2.0250 0.5550 ;
        RECT 1.7250 0.1500 1.8825 0.2550 ;
        RECT 1.4775 0.7800 1.8375 0.9000 ;
        RECT 1.4400 0.3300 1.7400 0.4050 ;
        RECT 1.5150 0.1500 1.6500 0.2550 ;
        RECT 1.2900 0.1500 1.5150 0.2325 ;
        RECT 1.3050 0.3075 1.4400 0.4050 ;
        RECT 1.3275 0.6300 1.4025 0.8325 ;
        RECT 1.1925 0.4800 1.2675 0.5850 ;
        RECT 1.0125 0.3825 1.1175 0.6825 ;
        RECT 0.8850 0.7950 1.0500 0.9000 ;
        RECT 0.8400 0.1575 1.0050 0.2775 ;
        RECT 0.8400 0.5100 0.9075 0.6600 ;
        RECT 0.6000 0.3525 0.9000 0.4275 ;
        RECT 0.6000 0.8250 0.8850 0.9000 ;
        RECT 0.6750 0.1575 0.8400 0.2625 ;
        RECT 0.7350 0.5100 0.8400 0.7350 ;
        RECT 0.5250 0.5025 0.6600 0.7500 ;
        RECT 0.5250 0.1800 0.6000 0.4275 ;
        RECT 0.3450 0.2550 0.4500 0.4500 ;
        RECT 0.3150 0.5250 0.4500 0.6900 ;
        RECT 0.1650 0.2550 0.3450 0.3300 ;
        RECT 0.2700 0.5250 0.3150 0.6150 ;
        RECT 0.1875 0.4725 0.2700 0.6150 ;
        RECT 0.1125 0.7050 0.1800 0.8850 ;
        RECT 0.1125 0.1950 0.1650 0.3300 ;
        RECT 0.0375 0.1950 0.1125 0.8850 ;
        LAYER VIA1 ;
        RECT 2.2500 0.2625 2.3250 0.3375 ;
        RECT 2.0475 0.8175 2.1225 0.8925 ;
        RECT 1.6875 0.8100 1.7625 0.8850 ;
        RECT 1.5300 0.1575 1.6050 0.2325 ;
        RECT 1.3725 0.3300 1.4475 0.4050 ;
        RECT 1.3275 0.7125 1.4025 0.7875 ;
        RECT 0.9300 0.8100 1.0050 0.8850 ;
        RECT 0.8850 0.2025 0.9600 0.2775 ;
        RECT 0.7425 0.6075 0.8175 0.6825 ;
        RECT 0.1050 0.7650 0.1800 0.8400 ;
        LAYER M2 ;
        RECT 2.0625 0.2625 2.3700 0.3375 ;
        RECT 2.0625 0.8175 2.1675 0.8925 ;
        RECT 1.9875 0.2625 2.0625 0.8925 ;
        RECT 1.6875 0.1575 1.7625 0.9375 ;
        RECT 0.9750 0.1575 1.6875 0.2325 ;
        RECT 1.0200 0.8625 1.6875 0.9375 ;
        RECT 1.5375 0.3300 1.6125 0.7875 ;
        RECT 1.3275 0.3300 1.5375 0.4050 ;
        RECT 1.2825 0.7125 1.5375 0.7875 ;
        RECT 0.9150 0.7650 1.0200 0.9375 ;
        RECT 0.8700 0.1575 0.9750 0.3225 ;
        RECT 0.8025 0.5625 0.8325 0.7275 ;
        RECT 0.7275 0.5625 0.8025 0.9375 ;
        RECT 0.1950 0.8625 0.7275 0.9375 ;
        RECT 0.0900 0.7200 0.1950 0.9375 ;
    END
END MUX3N_0011


MACRO MUX3N_0111
    CLASS CORE ;
    FOREIGN MUX3N_0111 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.7800 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 3.0975 0.2700 3.4125 0.7575 ;
        VIA 3.2550 0.3300 VIA12_slot ;
        VIA 3.2550 0.6975 VIA12_slot ;
        END
    END ZN
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.9125 0.1125 2.3775 0.1875 ;
        RECT 1.8375 0.1125 1.9125 0.6000 ;
        VIA 1.8750 0.5175 VIA12_square ;
        END
    END S1
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.4275 0.1125 0.7200 0.1875 ;
        RECT 0.4275 0.2625 0.6450 0.3375 ;
        RECT 0.3525 0.1125 0.4275 0.6900 ;
        RECT 0.1800 0.1125 0.3525 0.1875 ;
        VIA 0.5625 0.3000 VIA12_square ;
        VIA 0.3900 0.6075 VIA12_square ;
        END
    END S0
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 2.1975 0.5625 2.6625 0.6375 ;
        VIA 2.3250 0.6000 VIA12_square ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.9525 0.5625 1.4175 0.6375 ;
        VIA 1.0725 0.6000 VIA12_square ;
        END
    END I1
    PIN I0
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.6375 0.4125 1.1175 0.4875 ;
        RECT 0.5325 0.4125 0.6375 0.7500 ;
        VIA 0.5850 0.6675 VIA12_square ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 3.7125 -0.0750 3.7800 0.0750 ;
        RECT 3.6375 -0.0750 3.7125 0.3075 ;
        RECT 3.3150 -0.0750 3.6375 0.0750 ;
        RECT 3.1950 -0.0750 3.3150 0.2025 ;
        RECT 2.8950 -0.0750 3.1950 0.0750 ;
        RECT 2.7750 -0.0750 2.8950 0.1950 ;
        RECT 2.4750 -0.0750 2.7750 0.0750 ;
        RECT 2.3550 -0.0750 2.4750 0.1800 ;
        RECT 1.1850 -0.0750 2.3550 0.0750 ;
        RECT 1.0800 -0.0750 1.1850 0.2475 ;
        RECT 0.3750 -0.0750 1.0800 0.0750 ;
        RECT 0.2550 -0.0750 0.3750 0.1800 ;
        RECT 0.0000 -0.0750 0.2550 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 3.7275 0.9750 3.7800 1.1250 ;
        RECT 3.6225 0.6375 3.7275 1.1250 ;
        RECT 3.3150 0.9750 3.6225 1.1250 ;
        RECT 3.1950 0.8250 3.3150 1.1250 ;
        RECT 2.8950 0.9750 3.1950 1.1250 ;
        RECT 2.7750 0.8325 2.8950 1.1250 ;
        RECT 2.4750 0.9750 2.7750 1.1250 ;
        RECT 2.3550 0.7875 2.4750 1.1250 ;
        RECT 1.2000 0.9750 2.3550 1.1250 ;
        RECT 1.1250 0.7875 1.2000 1.1250 ;
        RECT 0.3750 0.9750 1.1250 1.1250 ;
        RECT 0.2550 0.7650 0.3750 1.1250 ;
        RECT 0.0000 0.9750 0.2550 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 3.6450 0.2175 3.7050 0.2775 ;
        RECT 3.6450 0.6675 3.7050 0.7275 ;
        RECT 3.6450 0.8325 3.7050 0.8925 ;
        RECT 3.5400 0.4800 3.6000 0.5400 ;
        RECT 3.4350 0.3000 3.4950 0.3600 ;
        RECT 3.4350 0.6675 3.4950 0.7275 ;
        RECT 3.3300 0.4800 3.3900 0.5400 ;
        RECT 3.2250 0.1350 3.2850 0.1950 ;
        RECT 3.2250 0.8325 3.2850 0.8925 ;
        RECT 3.1200 0.4800 3.1800 0.5400 ;
        RECT 3.0150 0.3000 3.0750 0.3600 ;
        RECT 3.0150 0.6675 3.0750 0.7275 ;
        RECT 2.9100 0.4800 2.9700 0.5400 ;
        RECT 2.8050 0.1350 2.8650 0.1950 ;
        RECT 2.8050 0.8400 2.8650 0.9000 ;
        RECT 2.7000 0.4800 2.7600 0.5400 ;
        RECT 2.5950 0.2850 2.6550 0.3450 ;
        RECT 2.5950 0.6750 2.6550 0.7350 ;
        RECT 2.4900 0.4800 2.5500 0.5400 ;
        RECT 2.3850 0.1200 2.4450 0.1800 ;
        RECT 2.3850 0.8175 2.4450 0.8775 ;
        RECT 2.2800 0.4500 2.3400 0.5100 ;
        RECT 2.0700 0.3975 2.1300 0.4575 ;
        RECT 2.0700 0.6375 2.1300 0.6975 ;
        RECT 1.9650 0.1650 2.0250 0.2250 ;
        RECT 1.9650 0.8100 2.0250 0.8700 ;
        RECT 1.8600 0.4875 1.9200 0.5475 ;
        RECT 1.7550 0.1650 1.8150 0.2250 ;
        RECT 1.7550 0.8175 1.8150 0.8775 ;
        RECT 1.6500 0.3375 1.7100 0.3975 ;
        RECT 1.5450 0.1650 1.6050 0.2250 ;
        RECT 1.3350 0.3075 1.3950 0.3675 ;
        RECT 1.3350 0.7350 1.3950 0.7950 ;
        RECT 1.2300 0.4875 1.2900 0.5475 ;
        RECT 1.1250 0.1575 1.1850 0.2175 ;
        RECT 1.1250 0.8175 1.1850 0.8775 ;
        RECT 1.0200 0.4650 1.0800 0.5250 ;
        RECT 0.8100 0.3600 0.8700 0.4200 ;
        RECT 0.8100 0.6000 0.8700 0.6600 ;
        RECT 0.7050 0.1725 0.7650 0.2325 ;
        RECT 0.7050 0.8325 0.7650 0.8925 ;
        RECT 0.6000 0.5700 0.6600 0.6300 ;
        RECT 0.3900 0.3600 0.4500 0.4200 ;
        RECT 0.3900 0.6000 0.4500 0.6600 ;
        RECT 0.2850 0.1200 0.3450 0.1800 ;
        RECT 0.2850 0.7950 0.3450 0.8550 ;
        RECT 0.1875 0.5025 0.2475 0.5625 ;
        RECT 0.0750 0.1950 0.1350 0.2550 ;
        RECT 0.0750 0.7725 0.1350 0.8325 ;
        LAYER M1 ;
        RECT 2.9100 0.4725 3.6300 0.5475 ;
        RECT 2.9850 0.2775 3.5250 0.3825 ;
        RECT 2.9850 0.6450 3.5250 0.7500 ;
        RECT 2.8350 0.2700 2.9100 0.7575 ;
        RECT 2.6925 0.2700 2.8350 0.3750 ;
        RECT 2.5725 0.6525 2.8350 0.7575 ;
        RECT 2.5125 0.4500 2.7600 0.5700 ;
        RECT 2.5875 0.2550 2.6925 0.3750 ;
        RECT 2.4375 0.2625 2.5125 0.5700 ;
        RECT 2.2800 0.2625 2.4375 0.3375 ;
        RECT 2.2725 0.4125 2.3625 0.6825 ;
        RECT 2.2050 0.1500 2.2800 0.3375 ;
        RECT 2.2050 0.4125 2.2725 0.5625 ;
        RECT 1.9125 0.7800 2.2275 0.9000 ;
        RECT 1.8825 0.1500 2.2050 0.2400 ;
        RECT 1.4025 0.6300 2.1675 0.7050 ;
        RECT 2.0250 0.3675 2.1300 0.5550 ;
        RECT 1.2675 0.4800 2.0250 0.5550 ;
        RECT 1.7250 0.1500 1.8825 0.2550 ;
        RECT 1.4775 0.7800 1.8375 0.9000 ;
        RECT 1.4400 0.3300 1.7400 0.4050 ;
        RECT 1.5150 0.1500 1.6500 0.2550 ;
        RECT 1.2900 0.1500 1.5150 0.2325 ;
        RECT 1.3050 0.3075 1.4400 0.4050 ;
        RECT 1.3275 0.6300 1.4025 0.8325 ;
        RECT 1.1925 0.4800 1.2675 0.5850 ;
        RECT 1.0125 0.3825 1.1175 0.6825 ;
        RECT 0.8850 0.7950 1.0500 0.9000 ;
        RECT 0.8400 0.1575 1.0050 0.2775 ;
        RECT 0.8400 0.5100 0.9075 0.6600 ;
        RECT 0.6000 0.3525 0.9000 0.4275 ;
        RECT 0.6000 0.8250 0.8850 0.9000 ;
        RECT 0.6750 0.1575 0.8400 0.2625 ;
        RECT 0.7350 0.5100 0.8400 0.7350 ;
        RECT 0.5250 0.5025 0.6600 0.7500 ;
        RECT 0.5250 0.1800 0.6000 0.4275 ;
        RECT 0.3450 0.2550 0.4500 0.4500 ;
        RECT 0.3150 0.5250 0.4500 0.6900 ;
        RECT 0.1650 0.2550 0.3450 0.3300 ;
        RECT 0.2700 0.5250 0.3150 0.6150 ;
        RECT 0.1875 0.4725 0.2700 0.6150 ;
        RECT 0.1125 0.7050 0.1800 0.8850 ;
        RECT 0.1125 0.1950 0.1650 0.3300 ;
        RECT 0.0375 0.1950 0.1125 0.8850 ;
        LAYER VIA1 ;
        RECT 2.2500 0.2625 2.3250 0.3375 ;
        RECT 2.0475 0.8175 2.1225 0.8925 ;
        RECT 1.6875 0.8100 1.7625 0.8850 ;
        RECT 1.5300 0.1575 1.6050 0.2325 ;
        RECT 1.3725 0.3300 1.4475 0.4050 ;
        RECT 1.3275 0.7125 1.4025 0.7875 ;
        RECT 0.9300 0.8100 1.0050 0.8850 ;
        RECT 0.8850 0.2025 0.9600 0.2775 ;
        RECT 0.7425 0.6075 0.8175 0.6825 ;
        RECT 0.1050 0.7650 0.1800 0.8400 ;
        LAYER M2 ;
        RECT 2.0625 0.2625 2.3700 0.3375 ;
        RECT 2.0625 0.8175 2.1675 0.8925 ;
        RECT 1.9875 0.2625 2.0625 0.8925 ;
        RECT 1.6875 0.1575 1.7625 0.9375 ;
        RECT 0.9750 0.1575 1.6875 0.2325 ;
        RECT 1.0200 0.8625 1.6875 0.9375 ;
        RECT 1.5375 0.3300 1.6125 0.7875 ;
        RECT 1.3275 0.3300 1.5375 0.4050 ;
        RECT 1.2825 0.7125 1.5375 0.7875 ;
        RECT 0.9150 0.7650 1.0200 0.9375 ;
        RECT 0.8700 0.1575 0.9750 0.3225 ;
        RECT 0.8025 0.5625 0.8325 0.7275 ;
        RECT 0.7275 0.5625 0.8025 0.9375 ;
        RECT 0.1950 0.8625 0.7275 0.9375 ;
        RECT 0.0900 0.7200 0.1950 0.9375 ;
    END
END MUX3N_0111


MACRO MUX3N_1000
    CLASS CORE ;
    FOREIGN MUX3N_1000 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.5200 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 2.0625 0.2625 2.4525 0.3375 ;
        RECT 2.0625 0.7875 2.1375 0.8925 ;
        RECT 1.9875 0.2625 2.0625 0.8925 ;
        VIA 2.2425 0.3000 VIA12_square ;
        VIA 2.0625 0.8400 VIA12_square ;
        END
    END ZN
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.9125 0.1125 2.3775 0.1875 ;
        RECT 1.8375 0.1125 1.9125 0.6000 ;
        VIA 1.8750 0.5175 VIA12_square ;
        END
    END S1
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.4275 0.1125 0.7200 0.1875 ;
        RECT 0.4275 0.2625 0.6450 0.3375 ;
        RECT 0.3525 0.1125 0.4275 0.6900 ;
        RECT 0.1800 0.1125 0.3525 0.1875 ;
        VIA 0.5625 0.3000 VIA12_square ;
        VIA 0.3900 0.6075 VIA12_square ;
        END
    END S0
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 2.3775 0.3675 2.4525 0.6825 ;
        RECT 2.2725 0.5625 2.3775 0.6825 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.9525 0.5625 1.4175 0.6375 ;
        VIA 1.0725 0.6000 VIA12_square ;
        END
    END I1
    PIN I0
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.6375 0.4125 1.1175 0.4875 ;
        RECT 0.5325 0.4125 0.6375 0.7500 ;
        VIA 0.5850 0.6675 VIA12_square ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 2.4750 -0.0750 2.5200 0.0750 ;
        RECT 2.3550 -0.0750 2.4750 0.2175 ;
        RECT 1.1850 -0.0750 2.3550 0.0750 ;
        RECT 1.0800 -0.0750 1.1850 0.2475 ;
        RECT 0.3750 -0.0750 1.0800 0.0750 ;
        RECT 0.2550 -0.0750 0.3750 0.1800 ;
        RECT 0.0000 -0.0750 0.2550 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 2.4750 0.9750 2.5200 1.1250 ;
        RECT 2.3550 0.7875 2.4750 1.1250 ;
        RECT 1.2000 0.9750 2.3550 1.1250 ;
        RECT 1.1250 0.7875 1.2000 1.1250 ;
        RECT 0.3750 0.9750 1.1250 1.1250 ;
        RECT 0.2550 0.7875 0.3750 1.1250 ;
        RECT 0.0000 0.9750 0.2550 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 2.3850 0.1575 2.4450 0.2175 ;
        RECT 2.3850 0.8175 2.4450 0.8775 ;
        RECT 2.2800 0.5925 2.3400 0.6525 ;
        RECT 2.0700 0.3975 2.1300 0.4575 ;
        RECT 2.0700 0.6375 2.1300 0.6975 ;
        RECT 1.9650 0.1575 2.0250 0.2175 ;
        RECT 1.9650 0.8100 2.0250 0.8700 ;
        RECT 1.8600 0.4875 1.9200 0.5475 ;
        RECT 1.7550 0.1575 1.8150 0.2175 ;
        RECT 1.7550 0.8175 1.8150 0.8775 ;
        RECT 1.6500 0.3375 1.7100 0.3975 ;
        RECT 1.5450 0.1575 1.6050 0.2175 ;
        RECT 1.3350 0.3075 1.3950 0.3675 ;
        RECT 1.3350 0.8175 1.3950 0.8775 ;
        RECT 1.2300 0.4875 1.2900 0.5475 ;
        RECT 1.1250 0.1575 1.1850 0.2175 ;
        RECT 1.1250 0.8175 1.1850 0.8775 ;
        RECT 1.0200 0.4650 1.0800 0.5250 ;
        RECT 0.8100 0.3600 0.8700 0.4200 ;
        RECT 0.8100 0.6000 0.8700 0.6600 ;
        RECT 0.7050 0.1725 0.7650 0.2325 ;
        RECT 0.7050 0.8325 0.7650 0.8925 ;
        RECT 0.6000 0.5700 0.6600 0.6300 ;
        RECT 0.3900 0.3600 0.4500 0.4200 ;
        RECT 0.3900 0.6000 0.4500 0.6600 ;
        RECT 0.2850 0.1200 0.3450 0.1800 ;
        RECT 0.2850 0.8175 0.3450 0.8775 ;
        RECT 0.1875 0.5025 0.2475 0.5625 ;
        RECT 0.0750 0.1575 0.1350 0.2175 ;
        RECT 0.0750 0.8175 0.1350 0.8775 ;
        LAYER M1 ;
        RECT 2.2050 0.1500 2.2800 0.3825 ;
        RECT 1.9125 0.7800 2.2275 0.9000 ;
        RECT 1.8825 0.1500 2.2050 0.2400 ;
        RECT 1.4175 0.6300 2.1600 0.7050 ;
        RECT 2.0250 0.3675 2.1300 0.5550 ;
        RECT 1.2675 0.4800 2.0250 0.5550 ;
        RECT 1.7250 0.1500 1.8825 0.2550 ;
        RECT 1.5000 0.7800 1.8375 0.9000 ;
        RECT 1.4400 0.3300 1.7400 0.4050 ;
        RECT 1.5150 0.1500 1.6500 0.2550 ;
        RECT 1.2900 0.1500 1.5150 0.2325 ;
        RECT 1.3050 0.3075 1.4400 0.4050 ;
        RECT 1.3425 0.6300 1.4175 0.9000 ;
        RECT 1.3125 0.7950 1.3425 0.9000 ;
        RECT 1.1925 0.4800 1.2675 0.5850 ;
        RECT 1.0125 0.3825 1.1175 0.6825 ;
        RECT 0.8850 0.7950 1.0500 0.9000 ;
        RECT 0.8400 0.1575 1.0050 0.2775 ;
        RECT 0.8400 0.5100 0.9075 0.6600 ;
        RECT 0.6000 0.3525 0.9000 0.4275 ;
        RECT 0.6000 0.8250 0.8850 0.9000 ;
        RECT 0.6750 0.1575 0.8400 0.2625 ;
        RECT 0.7350 0.5100 0.8400 0.7350 ;
        RECT 0.5250 0.5025 0.6600 0.7500 ;
        RECT 0.5250 0.1800 0.6000 0.4275 ;
        RECT 0.3450 0.2550 0.4500 0.4500 ;
        RECT 0.3150 0.5250 0.4500 0.6900 ;
        RECT 0.1650 0.2550 0.3450 0.3300 ;
        RECT 0.2700 0.5250 0.3150 0.6150 ;
        RECT 0.1875 0.4725 0.2700 0.6150 ;
        RECT 0.1125 0.7050 0.1800 0.8850 ;
        RECT 0.1125 0.1575 0.1650 0.3300 ;
        RECT 0.0375 0.1575 0.1125 0.8850 ;
        LAYER VIA1 ;
        RECT 1.6875 0.8100 1.7625 0.8850 ;
        RECT 1.5300 0.1575 1.6050 0.2325 ;
        RECT 1.3725 0.3300 1.4475 0.4050 ;
        RECT 1.3425 0.7125 1.4175 0.7875 ;
        RECT 0.9300 0.8100 1.0050 0.8850 ;
        RECT 0.8850 0.2025 0.9600 0.2775 ;
        RECT 0.7425 0.6075 0.8175 0.6825 ;
        RECT 0.1050 0.7650 0.1800 0.8400 ;
        LAYER M2 ;
        RECT 1.6875 0.1575 1.7625 0.9375 ;
        RECT 0.9750 0.1575 1.6875 0.2325 ;
        RECT 1.0200 0.8625 1.6875 0.9375 ;
        RECT 1.5375 0.3300 1.6125 0.7875 ;
        RECT 1.3275 0.3300 1.5375 0.4050 ;
        RECT 1.2825 0.7125 1.5375 0.7875 ;
        RECT 0.9150 0.7650 1.0200 0.9375 ;
        RECT 0.8700 0.1575 0.9750 0.3225 ;
        RECT 0.8025 0.5625 0.8325 0.7275 ;
        RECT 0.7275 0.5625 0.8025 0.9375 ;
        RECT 0.1950 0.8625 0.7275 0.9375 ;
        RECT 0.0900 0.7200 0.1950 0.9375 ;
    END
END MUX3N_1000


MACRO MUX3N_1010
    CLASS CORE ;
    FOREIGN MUX3N_1010 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.1500 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 3.0375 0.2175 3.1125 0.8325 ;
        RECT 3.0075 0.2175 3.0375 0.3825 ;
        RECT 3.0075 0.6675 3.0375 0.8325 ;
        END
    END ZN
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.9125 0.1125 2.3775 0.1875 ;
        RECT 1.8375 0.1125 1.9125 0.6000 ;
        VIA 1.8750 0.5175 VIA12_square ;
        END
    END S1
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.4275 0.1125 0.7200 0.1875 ;
        RECT 0.4275 0.2625 0.6450 0.3375 ;
        RECT 0.3525 0.1125 0.4275 0.6900 ;
        RECT 0.1800 0.1125 0.3525 0.1875 ;
        VIA 0.5625 0.3000 VIA12_square ;
        VIA 0.3900 0.6075 VIA12_square ;
        END
    END S0
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 2.1975 0.5625 2.6625 0.6375 ;
        VIA 2.3250 0.6000 VIA12_square ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.9525 0.5625 1.4175 0.6375 ;
        VIA 1.0725 0.6000 VIA12_square ;
        END
    END I1
    PIN I0
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.6375 0.4125 1.1175 0.4875 ;
        RECT 0.5325 0.4125 0.6375 0.7500 ;
        VIA 0.5850 0.6675 VIA12_square ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 2.8875 -0.0750 3.1500 0.0750 ;
        RECT 2.7825 -0.0750 2.8875 0.2925 ;
        RECT 2.4750 -0.0750 2.7825 0.0750 ;
        RECT 2.3550 -0.0750 2.4750 0.1800 ;
        RECT 1.1850 -0.0750 2.3550 0.0750 ;
        RECT 1.0800 -0.0750 1.1850 0.2475 ;
        RECT 0.3750 -0.0750 1.0800 0.0750 ;
        RECT 0.2550 -0.0750 0.3750 0.1800 ;
        RECT 0.0000 -0.0750 0.2550 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 2.8875 0.9750 3.1500 1.1250 ;
        RECT 2.7825 0.6375 2.8875 1.1250 ;
        RECT 2.4750 0.9750 2.7825 1.1250 ;
        RECT 2.3550 0.7875 2.4750 1.1250 ;
        RECT 1.2000 0.9750 2.3550 1.1250 ;
        RECT 1.1250 0.7875 1.2000 1.1250 ;
        RECT 0.3750 0.9750 1.1250 1.1250 ;
        RECT 0.2550 0.7650 0.3750 1.1250 ;
        RECT 0.0000 0.9750 0.2550 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 3.0150 0.2700 3.0750 0.3300 ;
        RECT 3.0150 0.7200 3.0750 0.7800 ;
        RECT 2.9025 0.4725 2.9625 0.5325 ;
        RECT 2.8050 0.2100 2.8650 0.2700 ;
        RECT 2.8050 0.6675 2.8650 0.7275 ;
        RECT 2.8050 0.8325 2.8650 0.8925 ;
        RECT 2.5950 0.2700 2.6550 0.3300 ;
        RECT 2.5950 0.7500 2.6550 0.8100 ;
        RECT 2.4825 0.4800 2.5425 0.5400 ;
        RECT 2.3850 0.1200 2.4450 0.1800 ;
        RECT 2.3850 0.8175 2.4450 0.8775 ;
        RECT 2.2800 0.4500 2.3400 0.5100 ;
        RECT 2.0700 0.3975 2.1300 0.4575 ;
        RECT 2.0700 0.6375 2.1300 0.6975 ;
        RECT 1.9650 0.1650 2.0250 0.2250 ;
        RECT 1.9650 0.8100 2.0250 0.8700 ;
        RECT 1.8600 0.4875 1.9200 0.5475 ;
        RECT 1.7550 0.1650 1.8150 0.2250 ;
        RECT 1.7550 0.8175 1.8150 0.8775 ;
        RECT 1.6500 0.3375 1.7100 0.3975 ;
        RECT 1.5450 0.1650 1.6050 0.2250 ;
        RECT 1.3350 0.3075 1.3950 0.3675 ;
        RECT 1.3350 0.7350 1.3950 0.7950 ;
        RECT 1.2300 0.4875 1.2900 0.5475 ;
        RECT 1.1250 0.1575 1.1850 0.2175 ;
        RECT 1.1250 0.8175 1.1850 0.8775 ;
        RECT 1.0200 0.4650 1.0800 0.5250 ;
        RECT 0.8100 0.3600 0.8700 0.4200 ;
        RECT 0.8100 0.6000 0.8700 0.6600 ;
        RECT 0.7050 0.1725 0.7650 0.2325 ;
        RECT 0.7050 0.8325 0.7650 0.8925 ;
        RECT 0.6000 0.5700 0.6600 0.6300 ;
        RECT 0.3900 0.3600 0.4500 0.4200 ;
        RECT 0.3900 0.6000 0.4500 0.6600 ;
        RECT 0.2850 0.1200 0.3450 0.1800 ;
        RECT 0.2850 0.7950 0.3450 0.8550 ;
        RECT 0.1875 0.5025 0.2475 0.5625 ;
        RECT 0.0750 0.1950 0.1350 0.2550 ;
        RECT 0.0750 0.7725 0.1350 0.8325 ;
        LAYER M1 ;
        RECT 2.6925 0.4425 2.9625 0.5625 ;
        RECT 2.6175 0.2175 2.6925 0.8400 ;
        RECT 2.5875 0.2175 2.6175 0.3825 ;
        RECT 2.5875 0.7200 2.6175 0.8400 ;
        RECT 2.5125 0.4500 2.5425 0.5700 ;
        RECT 2.4375 0.2625 2.5125 0.5700 ;
        RECT 2.2800 0.2625 2.4375 0.3375 ;
        RECT 2.2725 0.4125 2.3625 0.6825 ;
        RECT 2.2050 0.1500 2.2800 0.3375 ;
        RECT 2.2050 0.4125 2.2725 0.5625 ;
        RECT 1.9125 0.7800 2.2275 0.9000 ;
        RECT 1.8825 0.1500 2.2050 0.2400 ;
        RECT 1.4025 0.6300 2.1675 0.7050 ;
        RECT 2.0250 0.3675 2.1300 0.5550 ;
        RECT 1.2675 0.4800 2.0250 0.5550 ;
        RECT 1.7250 0.1500 1.8825 0.2550 ;
        RECT 1.4775 0.7800 1.8375 0.9000 ;
        RECT 1.4400 0.3300 1.7400 0.4050 ;
        RECT 1.5150 0.1500 1.6500 0.2550 ;
        RECT 1.2900 0.1500 1.5150 0.2325 ;
        RECT 1.3050 0.3075 1.4400 0.4050 ;
        RECT 1.3275 0.6300 1.4025 0.8325 ;
        RECT 1.1925 0.4800 1.2675 0.5850 ;
        RECT 1.0125 0.3825 1.1175 0.6825 ;
        RECT 0.8850 0.7950 1.0500 0.9000 ;
        RECT 0.8400 0.1575 1.0050 0.2775 ;
        RECT 0.8400 0.5100 0.9075 0.6600 ;
        RECT 0.6000 0.3525 0.9000 0.4275 ;
        RECT 0.6000 0.8250 0.8850 0.9000 ;
        RECT 0.6750 0.1575 0.8400 0.2625 ;
        RECT 0.7350 0.5100 0.8400 0.7350 ;
        RECT 0.5250 0.5025 0.6600 0.7500 ;
        RECT 0.5250 0.1800 0.6000 0.4275 ;
        RECT 0.3450 0.2550 0.4500 0.4500 ;
        RECT 0.3150 0.5250 0.4500 0.6900 ;
        RECT 0.1650 0.2550 0.3450 0.3300 ;
        RECT 0.2700 0.5250 0.3150 0.6150 ;
        RECT 0.1875 0.4725 0.2700 0.6150 ;
        RECT 0.1125 0.7050 0.1800 0.8850 ;
        RECT 0.1125 0.1950 0.1650 0.3300 ;
        RECT 0.0375 0.1950 0.1125 0.8850 ;
        LAYER VIA1 ;
        RECT 2.2500 0.2625 2.3250 0.3375 ;
        RECT 2.0475 0.8175 2.1225 0.8925 ;
        RECT 1.6875 0.8100 1.7625 0.8850 ;
        RECT 1.5300 0.1575 1.6050 0.2325 ;
        RECT 1.3725 0.3300 1.4475 0.4050 ;
        RECT 1.3275 0.7125 1.4025 0.7875 ;
        RECT 0.9300 0.8100 1.0050 0.8850 ;
        RECT 0.8850 0.2025 0.9600 0.2775 ;
        RECT 0.7425 0.6075 0.8175 0.6825 ;
        RECT 0.1050 0.7650 0.1800 0.8400 ;
        LAYER M2 ;
        RECT 2.0625 0.2625 2.3700 0.3375 ;
        RECT 2.0625 0.8175 2.1675 0.8925 ;
        RECT 1.9875 0.2625 2.0625 0.8925 ;
        RECT 1.6875 0.1575 1.7625 0.9375 ;
        RECT 0.9750 0.1575 1.6875 0.2325 ;
        RECT 1.0200 0.8625 1.6875 0.9375 ;
        RECT 1.5375 0.3300 1.6125 0.7875 ;
        RECT 1.3275 0.3300 1.5375 0.4050 ;
        RECT 1.2825 0.7125 1.5375 0.7875 ;
        RECT 0.9150 0.7650 1.0200 0.9375 ;
        RECT 0.8700 0.1575 0.9750 0.3225 ;
        RECT 0.8025 0.5625 0.8325 0.7275 ;
        RECT 0.7275 0.5625 0.8025 0.9375 ;
        RECT 0.1950 0.8625 0.7275 0.9375 ;
        RECT 0.0900 0.7200 0.1950 0.9375 ;
    END
END MUX3N_1010


MACRO MUX3_0111
    CLASS CORE ;
    FOREIGN MUX3_0111 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.8300 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 4.1475 0.2700 4.4625 0.7575 ;
        VIA 4.3050 0.3300 VIA12_slot ;
        VIA 4.3050 0.6975 VIA12_slot ;
        END
    END Z
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 2.8725 0.5625 3.3375 0.6375 ;
        RECT 2.7975 0.4050 2.8725 0.6375 ;
        VIA 2.8350 0.4875 VIA12_square ;
        END
    END S1
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.2450 0.3525 1.4175 0.4575 ;
        RECT 1.1700 0.1125 1.2450 0.4575 ;
        RECT 0.4275 0.1125 1.1700 0.1875 ;
        RECT 0.3525 0.1125 0.4275 0.6450 ;
        VIA 1.3425 0.4050 VIA12_square ;
        VIA 0.3900 0.5625 VIA12_square ;
        END
    END S0
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 3.6225 0.4125 3.7275 0.5850 ;
        RECT 3.1575 0.4125 3.6225 0.4875 ;
        VIA 3.6750 0.5100 VIA12_square ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.7325 0.4125 2.1975 0.4875 ;
        VIA 2.1075 0.4500 VIA12_square ;
        END
    END I1
    PIN I0
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.0125 0.2625 1.0875 0.6075 ;
        RECT 0.5475 0.2625 1.0125 0.3375 ;
        VIA 1.0500 0.5250 VIA12_square ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 4.7625 -0.0750 4.8300 0.0750 ;
        RECT 4.6875 -0.0750 4.7625 0.3075 ;
        RECT 4.3650 -0.0750 4.6875 0.0750 ;
        RECT 4.2450 -0.0750 4.3650 0.2025 ;
        RECT 3.9225 -0.0750 4.2450 0.0750 ;
        RECT 3.8475 -0.0750 3.9225 0.3075 ;
        RECT 3.5250 -0.0750 3.8475 0.0750 ;
        RECT 3.4050 -0.0750 3.5250 0.2250 ;
        RECT 2.2350 -0.0750 3.4050 0.0750 ;
        RECT 2.1600 -0.0750 2.2350 0.2475 ;
        RECT 1.8450 -0.0750 2.1600 0.0750 ;
        RECT 1.7250 -0.0750 1.8450 0.2250 ;
        RECT 0.7950 -0.0750 1.7250 0.0750 ;
        RECT 0.6750 -0.0750 0.7950 0.2175 ;
        RECT 0.3675 -0.0750 0.6750 0.0750 ;
        RECT 0.2625 -0.0750 0.3675 0.2400 ;
        RECT 0.0000 -0.0750 0.2625 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 4.7775 0.9750 4.8300 1.1250 ;
        RECT 4.6725 0.6375 4.7775 1.1250 ;
        RECT 4.3650 0.9750 4.6725 1.1250 ;
        RECT 4.2450 0.8250 4.3650 1.1250 ;
        RECT 3.9375 0.9750 4.2450 1.1250 ;
        RECT 3.8325 0.6675 3.9375 1.1250 ;
        RECT 3.5400 0.9750 3.8325 1.1250 ;
        RECT 3.4350 0.8025 3.5400 1.1250 ;
        RECT 2.2425 0.9750 3.4350 1.1250 ;
        RECT 2.1675 0.7650 2.2425 1.1250 ;
        RECT 1.8375 0.9750 2.1675 1.1250 ;
        RECT 1.7325 0.7800 1.8375 1.1250 ;
        RECT 0.7950 0.9750 1.7325 1.1250 ;
        RECT 0.6750 0.8325 0.7950 1.1250 ;
        RECT 0.3600 0.9750 0.6750 1.1250 ;
        RECT 0.2700 0.7950 0.3600 1.1250 ;
        RECT 0.0000 0.9750 0.2700 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 4.6950 0.2175 4.7550 0.2775 ;
        RECT 4.6950 0.6675 4.7550 0.7275 ;
        RECT 4.6950 0.8325 4.7550 0.8925 ;
        RECT 4.5900 0.4800 4.6500 0.5400 ;
        RECT 4.4850 0.3000 4.5450 0.3600 ;
        RECT 4.4850 0.6675 4.5450 0.7275 ;
        RECT 4.3800 0.4800 4.4400 0.5400 ;
        RECT 4.2750 0.1350 4.3350 0.1950 ;
        RECT 4.2750 0.8325 4.3350 0.8925 ;
        RECT 4.1700 0.4800 4.2300 0.5400 ;
        RECT 4.0650 0.3000 4.1250 0.3600 ;
        RECT 4.0650 0.6675 4.1250 0.7275 ;
        RECT 3.9600 0.4800 4.0200 0.5400 ;
        RECT 3.8550 0.2175 3.9150 0.2775 ;
        RECT 3.8550 0.6900 3.9150 0.7500 ;
        RECT 3.8550 0.8550 3.9150 0.9150 ;
        RECT 3.7500 0.4800 3.8100 0.5400 ;
        RECT 3.6450 0.2775 3.7050 0.3375 ;
        RECT 3.6450 0.6900 3.7050 0.7500 ;
        RECT 3.5400 0.4800 3.6000 0.5400 ;
        RECT 3.4350 0.1575 3.4950 0.2175 ;
        RECT 3.4350 0.8325 3.4950 0.8925 ;
        RECT 3.2250 0.1800 3.2850 0.2400 ;
        RECT 3.2250 0.8100 3.2850 0.8700 ;
        RECT 3.1200 0.3750 3.1800 0.4350 ;
        RECT 3.1200 0.6150 3.1800 0.6750 ;
        RECT 3.0150 0.1725 3.0750 0.2325 ;
        RECT 3.0150 0.8100 3.0750 0.8700 ;
        RECT 2.9100 0.4575 2.9700 0.5175 ;
        RECT 2.8050 0.1800 2.8650 0.2400 ;
        RECT 2.8050 0.8100 2.8650 0.8700 ;
        RECT 2.7000 0.6225 2.7600 0.6825 ;
        RECT 2.5950 0.1650 2.6550 0.2250 ;
        RECT 2.3850 0.3075 2.4450 0.3675 ;
        RECT 2.3850 0.7050 2.4450 0.7650 ;
        RECT 2.2800 0.4800 2.3400 0.5400 ;
        RECT 2.1750 0.1575 2.2350 0.2175 ;
        RECT 2.1750 0.7950 2.2350 0.8550 ;
        RECT 2.0700 0.4725 2.1300 0.5325 ;
        RECT 1.9650 0.1650 2.0250 0.2250 ;
        RECT 1.9650 0.6600 2.0250 0.7200 ;
        RECT 1.8600 0.4725 1.9200 0.5325 ;
        RECT 1.7550 0.1575 1.8150 0.2175 ;
        RECT 1.7550 0.8025 1.8150 0.8625 ;
        RECT 1.5450 0.1800 1.6050 0.2400 ;
        RECT 1.5450 0.8100 1.6050 0.8700 ;
        RECT 1.4400 0.3600 1.5000 0.4200 ;
        RECT 1.4400 0.6000 1.5000 0.6600 ;
        RECT 1.3350 0.1650 1.3950 0.2250 ;
        RECT 1.3350 0.8175 1.3950 0.8775 ;
        RECT 1.1250 0.1725 1.1850 0.2325 ;
        RECT 1.1250 0.8175 1.1850 0.8775 ;
        RECT 1.0200 0.4950 1.0800 0.5550 ;
        RECT 0.9150 0.2025 0.9750 0.2625 ;
        RECT 0.9150 0.6900 0.9750 0.7500 ;
        RECT 0.8100 0.5100 0.8700 0.5700 ;
        RECT 0.7050 0.1575 0.7650 0.2175 ;
        RECT 0.7050 0.8325 0.7650 0.8925 ;
        RECT 0.6000 0.5100 0.6600 0.5700 ;
        RECT 0.4950 0.1725 0.5550 0.2325 ;
        RECT 0.4950 0.7875 0.5550 0.8475 ;
        RECT 0.3900 0.3600 0.4500 0.4200 ;
        RECT 0.3900 0.6000 0.4500 0.6600 ;
        RECT 0.2850 0.1575 0.3450 0.2175 ;
        RECT 0.2850 0.8250 0.3450 0.8850 ;
        RECT 0.1875 0.5550 0.2475 0.6150 ;
        RECT 0.0750 0.2025 0.1350 0.2625 ;
        RECT 0.0750 0.7725 0.1350 0.8325 ;
        LAYER M1 ;
        RECT 3.9075 0.4575 4.6725 0.5625 ;
        RECT 4.0350 0.2775 4.5750 0.3825 ;
        RECT 4.0350 0.6450 4.5750 0.7500 ;
        RECT 3.5175 0.4575 3.8325 0.5625 ;
        RECT 3.6375 0.2475 3.7125 0.3750 ;
        RECT 3.6375 0.6525 3.7125 0.7800 ;
        RECT 3.3300 0.3000 3.6375 0.3750 ;
        RECT 3.3600 0.6525 3.6375 0.7275 ;
        RECT 3.2850 0.6525 3.3600 0.9000 ;
        RECT 3.2550 0.1500 3.3300 0.3750 ;
        RECT 3.2250 0.7800 3.2850 0.9000 ;
        RECT 3.2250 0.1500 3.2550 0.2700 ;
        RECT 3.0975 0.5700 3.2100 0.6750 ;
        RECT 3.0750 0.3450 3.1800 0.4650 ;
        RECT 2.8050 0.1500 3.1500 0.2700 ;
        RECT 2.9400 0.7500 3.1500 0.9000 ;
        RECT 2.8950 0.6000 3.0975 0.6750 ;
        RECT 3.0000 0.3900 3.0750 0.4650 ;
        RECT 2.9250 0.3900 3.0000 0.5250 ;
        RECT 2.7750 0.4500 2.9250 0.5250 ;
        RECT 2.8200 0.6000 2.8950 0.6900 ;
        RECT 2.5275 0.7800 2.8650 0.9000 ;
        RECT 2.4525 0.6150 2.8200 0.6900 ;
        RECT 2.7000 0.4500 2.7750 0.5400 ;
        RECT 2.3400 0.1500 2.7000 0.2325 ;
        RECT 2.3175 0.4650 2.7000 0.5400 ;
        RECT 2.3250 0.3075 2.6550 0.3900 ;
        RECT 2.3775 0.6150 2.4525 0.8100 ;
        RECT 2.2425 0.4650 2.3175 0.5700 ;
        RECT 2.0700 0.3675 2.1675 0.5550 ;
        RECT 1.8375 0.4500 2.0700 0.5550 ;
        RECT 1.9950 0.1500 2.0550 0.2400 ;
        RECT 1.9575 0.6300 2.0325 0.7500 ;
        RECT 1.9200 0.1500 1.9950 0.3750 ;
        RECT 1.6575 0.6300 1.9575 0.7050 ;
        RECT 1.6500 0.3000 1.9200 0.3750 ;
        RECT 1.5825 0.6300 1.6575 0.9000 ;
        RECT 1.5750 0.1500 1.6500 0.3750 ;
        RECT 1.5450 0.7800 1.5825 0.9000 ;
        RECT 1.5450 0.1500 1.5750 0.2700 ;
        RECT 1.2900 0.5550 1.5075 0.7050 ;
        RECT 1.2900 0.3300 1.5000 0.4800 ;
        RECT 1.1025 0.1500 1.4700 0.2550 ;
        RECT 1.1025 0.7950 1.4700 0.9000 ;
        RECT 1.0125 0.4425 1.2150 0.6075 ;
        RECT 0.6000 0.6825 1.0050 0.7575 ;
        RECT 0.9075 0.1725 0.9825 0.3675 ;
        RECT 0.7425 0.4425 0.9375 0.6075 ;
        RECT 0.6000 0.2925 0.9075 0.3675 ;
        RECT 0.5925 0.4800 0.6675 0.6000 ;
        RECT 0.5250 0.1500 0.6000 0.3675 ;
        RECT 0.5250 0.6825 0.6000 0.8775 ;
        RECT 0.4500 0.5250 0.5925 0.6000 ;
        RECT 0.4725 0.1500 0.5250 0.2550 ;
        RECT 0.4875 0.7575 0.5250 0.8775 ;
        RECT 0.1575 0.3300 0.4500 0.4500 ;
        RECT 0.3450 0.5250 0.4500 0.6900 ;
        RECT 0.1875 0.5250 0.3450 0.6450 ;
        RECT 0.1125 0.7275 0.1950 0.9000 ;
        RECT 0.1125 0.1725 0.1575 0.4500 ;
        RECT 0.0375 0.1725 0.1125 0.9000 ;
        LAYER VIA1 ;
        RECT 3.9450 0.4725 4.0200 0.5475 ;
        RECT 3.0375 0.1650 3.1125 0.2400 ;
        RECT 3.0075 0.7650 3.0825 0.8400 ;
        RECT 2.5650 0.8100 2.6400 0.8850 ;
        RECT 2.5425 0.6150 2.6175 0.6900 ;
        RECT 2.5350 0.3150 2.6100 0.3900 ;
        RECT 2.3850 0.1575 2.4600 0.2325 ;
        RECT 1.3575 0.1650 1.4325 0.2400 ;
        RECT 1.3575 0.8100 1.4325 0.8850 ;
        RECT 1.3050 0.5925 1.3800 0.6675 ;
        RECT 0.7425 0.4875 0.8175 0.5625 ;
        RECT 0.1050 0.7725 0.1800 0.8475 ;
        LAYER M2 ;
        RECT 3.8925 0.4575 4.0575 0.5625 ;
        RECT 3.8175 0.2625 3.8925 0.7875 ;
        RECT 3.1500 0.2625 3.8175 0.3375 ;
        RECT 3.0975 0.7125 3.8175 0.7875 ;
        RECT 2.9925 0.1500 3.1500 0.3375 ;
        RECT 2.9925 0.7125 3.0975 0.8775 ;
        RECT 2.5275 0.7950 2.6775 0.9000 ;
        RECT 2.5875 0.3150 2.6625 0.6900 ;
        RECT 2.4900 0.3150 2.5875 0.3900 ;
        RECT 2.4975 0.6150 2.5875 0.6900 ;
        RECT 1.6125 0.8100 2.5275 0.8850 ;
        RECT 2.3400 0.1500 2.5050 0.2400 ;
        RECT 1.6125 0.1650 2.3400 0.2400 ;
        RECT 1.5375 0.1650 1.6125 0.8850 ;
        RECT 1.4700 0.1650 1.5375 0.2550 ;
        RECT 1.4700 0.7950 1.5375 0.8850 ;
        RECT 1.3200 0.1500 1.4700 0.2550 ;
        RECT 1.3200 0.7950 1.4700 0.9000 ;
        RECT 1.2450 0.5775 1.4175 0.6825 ;
        RECT 1.1700 0.5775 1.2450 0.8850 ;
        RECT 0.8175 0.8100 1.1700 0.8850 ;
        RECT 0.7425 0.4425 0.8175 0.8850 ;
        RECT 0.1950 0.8100 0.7425 0.8850 ;
        RECT 0.0900 0.7350 0.1950 0.8850 ;
    END
END MUX3_0111


MACRO MUX3_1010
    CLASS CORE ;
    FOREIGN MUX3_1010 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.7300 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 2.6175 0.2175 2.6925 0.8325 ;
        RECT 2.5875 0.2175 2.6175 0.3825 ;
        RECT 2.5875 0.6675 2.6175 0.8325 ;
        END
    END Z
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.9125 0.1125 2.3775 0.1875 ;
        RECT 1.8375 0.1125 1.9125 0.6000 ;
        VIA 1.8750 0.5175 VIA12_square ;
        END
    END S1
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.4275 0.1125 0.7200 0.1875 ;
        RECT 0.4275 0.2625 0.6450 0.3375 ;
        RECT 0.3525 0.1125 0.4275 0.6900 ;
        RECT 0.1800 0.1125 0.3525 0.1875 ;
        VIA 0.5625 0.3000 VIA12_square ;
        VIA 0.3900 0.6075 VIA12_square ;
        END
    END S0
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 2.1975 0.5625 2.6625 0.6375 ;
        VIA 2.3250 0.6000 VIA12_square ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.9525 0.5625 1.4175 0.6375 ;
        VIA 1.0725 0.6000 VIA12_square ;
        END
    END I1
    PIN I0
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.6375 0.4125 1.1175 0.4875 ;
        RECT 0.5325 0.4125 0.6375 0.7500 ;
        VIA 0.5850 0.6675 VIA12_square ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 2.4750 -0.0750 2.7300 0.0750 ;
        RECT 2.3550 -0.0750 2.4750 0.1800 ;
        RECT 1.1850 -0.0750 2.3550 0.0750 ;
        RECT 1.0800 -0.0750 1.1850 0.2475 ;
        RECT 0.3750 -0.0750 1.0800 0.0750 ;
        RECT 0.2550 -0.0750 0.3750 0.1800 ;
        RECT 0.0000 -0.0750 0.2550 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 2.4750 0.9750 2.7300 1.1250 ;
        RECT 2.3550 0.7950 2.4750 1.1250 ;
        RECT 1.2000 0.9750 2.3550 1.1250 ;
        RECT 1.1250 0.7950 1.2000 1.1250 ;
        RECT 0.3750 0.9750 1.1250 1.1250 ;
        RECT 0.2550 0.7650 0.3750 1.1250 ;
        RECT 0.0000 0.9750 0.2550 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 2.5950 0.2700 2.6550 0.3300 ;
        RECT 2.5950 0.7200 2.6550 0.7800 ;
        RECT 2.4825 0.4800 2.5425 0.5400 ;
        RECT 2.3850 0.1200 2.4450 0.1800 ;
        RECT 2.3850 0.8250 2.4450 0.8850 ;
        RECT 2.2800 0.4500 2.3400 0.5100 ;
        RECT 2.0700 0.3975 2.1300 0.4575 ;
        RECT 2.0700 0.6375 2.1300 0.6975 ;
        RECT 1.9650 0.1650 2.0250 0.2250 ;
        RECT 1.9650 0.8100 2.0250 0.8700 ;
        RECT 1.8600 0.4875 1.9200 0.5475 ;
        RECT 1.7550 0.1650 1.8150 0.2250 ;
        RECT 1.7550 0.8175 1.8150 0.8775 ;
        RECT 1.6500 0.3375 1.7100 0.3975 ;
        RECT 1.5450 0.1650 1.6050 0.2250 ;
        RECT 1.3350 0.3075 1.3950 0.3675 ;
        RECT 1.3350 0.7350 1.3950 0.7950 ;
        RECT 1.2300 0.4875 1.2900 0.5475 ;
        RECT 1.1250 0.1575 1.1850 0.2175 ;
        RECT 1.1250 0.8250 1.1850 0.8850 ;
        RECT 1.0200 0.4650 1.0800 0.5250 ;
        RECT 0.8100 0.3600 0.8700 0.4200 ;
        RECT 0.8100 0.6000 0.8700 0.6600 ;
        RECT 0.7050 0.1725 0.7650 0.2325 ;
        RECT 0.7050 0.8325 0.7650 0.8925 ;
        RECT 0.6000 0.5700 0.6600 0.6300 ;
        RECT 0.3900 0.3600 0.4500 0.4200 ;
        RECT 0.3900 0.6000 0.4500 0.6600 ;
        RECT 0.2850 0.1200 0.3450 0.1800 ;
        RECT 0.2850 0.7875 0.3450 0.8475 ;
        RECT 0.1875 0.5025 0.2475 0.5625 ;
        RECT 0.0750 0.2025 0.1350 0.2625 ;
        RECT 0.0750 0.7725 0.1350 0.8325 ;
        LAYER M1 ;
        RECT 2.5125 0.4500 2.5425 0.5700 ;
        RECT 2.4375 0.2625 2.5125 0.5700 ;
        RECT 2.2800 0.2625 2.4375 0.3375 ;
        RECT 2.2725 0.4125 2.3625 0.6825 ;
        RECT 2.2050 0.1500 2.2800 0.3375 ;
        RECT 2.2050 0.4125 2.2725 0.5625 ;
        RECT 1.9125 0.7800 2.2275 0.9000 ;
        RECT 1.8825 0.1500 2.2050 0.2400 ;
        RECT 1.4025 0.6300 2.1675 0.7050 ;
        RECT 2.0250 0.3675 2.1300 0.5550 ;
        RECT 1.2675 0.4800 2.0250 0.5550 ;
        RECT 1.7250 0.1500 1.8825 0.2550 ;
        RECT 1.4775 0.7800 1.8375 0.9000 ;
        RECT 1.4400 0.3300 1.7400 0.4050 ;
        RECT 1.5150 0.1500 1.6500 0.2550 ;
        RECT 1.2900 0.1500 1.5150 0.2325 ;
        RECT 1.3050 0.3075 1.4400 0.4050 ;
        RECT 1.3275 0.6300 1.4025 0.8325 ;
        RECT 1.1925 0.4800 1.2675 0.5850 ;
        RECT 1.0125 0.3825 1.1175 0.6825 ;
        RECT 0.8850 0.7950 1.0500 0.9000 ;
        RECT 0.8400 0.1575 1.0050 0.2775 ;
        RECT 0.8400 0.5100 0.9075 0.6600 ;
        RECT 0.6000 0.3525 0.9000 0.4275 ;
        RECT 0.6000 0.8250 0.8850 0.9000 ;
        RECT 0.6750 0.1575 0.8400 0.2625 ;
        RECT 0.7350 0.5100 0.8400 0.7350 ;
        RECT 0.5250 0.5025 0.6600 0.7500 ;
        RECT 0.5250 0.1800 0.6000 0.4275 ;
        RECT 0.3450 0.2550 0.4500 0.4500 ;
        RECT 0.3150 0.5250 0.4500 0.6900 ;
        RECT 0.1650 0.2550 0.3450 0.3300 ;
        RECT 0.2700 0.5250 0.3150 0.6150 ;
        RECT 0.1875 0.4725 0.2700 0.6150 ;
        RECT 0.1125 0.7050 0.1800 0.8850 ;
        RECT 0.1125 0.1725 0.1650 0.3300 ;
        RECT 0.0375 0.1725 0.1125 0.8850 ;
        LAYER VIA1 ;
        RECT 2.2500 0.2625 2.3250 0.3375 ;
        RECT 2.0475 0.8175 2.1225 0.8925 ;
        RECT 1.6875 0.8100 1.7625 0.8850 ;
        RECT 1.5300 0.1575 1.6050 0.2325 ;
        RECT 1.3725 0.3300 1.4475 0.4050 ;
        RECT 1.3275 0.7125 1.4025 0.7875 ;
        RECT 0.9300 0.8100 1.0050 0.8850 ;
        RECT 0.8850 0.2025 0.9600 0.2775 ;
        RECT 0.7425 0.6075 0.8175 0.6825 ;
        RECT 0.1050 0.7650 0.1800 0.8400 ;
        LAYER M2 ;
        RECT 2.0625 0.2625 2.3700 0.3375 ;
        RECT 2.0625 0.8175 2.1675 0.8925 ;
        RECT 1.9875 0.2625 2.0625 0.8925 ;
        RECT 1.6875 0.1575 1.7625 0.9375 ;
        RECT 0.9750 0.1575 1.6875 0.2325 ;
        RECT 1.0200 0.8625 1.6875 0.9375 ;
        RECT 1.5375 0.3300 1.6125 0.7875 ;
        RECT 1.3275 0.3300 1.5375 0.4050 ;
        RECT 1.2825 0.7125 1.5375 0.7875 ;
        RECT 0.9150 0.7650 1.0200 0.9375 ;
        RECT 0.8700 0.1575 0.9750 0.3225 ;
        RECT 0.8025 0.5625 0.8325 0.7275 ;
        RECT 0.7275 0.5625 0.8025 0.9375 ;
        RECT 0.1950 0.8625 0.7275 0.9375 ;
        RECT 0.0900 0.7200 0.1950 0.9375 ;
    END
END MUX3_1010


MACRO MUX4_1010
    CLASS CORE ;
    FOREIGN MUX4_1010 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.9900 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 3.0675 0.1125 3.6375 0.1875 ;
        RECT 3.0675 0.4800 3.2025 0.5550 ;
        RECT 2.9925 0.1125 3.0675 0.5550 ;
        VIA 3.1200 0.5175 VIA12_square ;
        END
    END S1
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.8450 0.1125 1.9200 0.4875 ;
        RECT 0.3225 0.1125 1.8450 0.1875 ;
        RECT 1.5300 0.4125 1.8450 0.4875 ;
        RECT 1.4550 0.4125 1.5300 0.7875 ;
        RECT 0.6450 0.7125 1.4550 0.7875 ;
        RECT 0.2175 0.1125 0.3225 0.3000 ;
        VIA 1.8825 0.3675 VIA12_square ;
        VIA 1.4925 0.6975 VIA12_square ;
        VIA 0.7575 0.7500 VIA12_square ;
        VIA 0.2700 0.2250 VIA12_square ;
        END
    END S0
    PIN I3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1425 0.5550 0.2550 0.6825 ;
        RECT 0.0675 0.3675 0.1425 0.6825 ;
        END
    END I3
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.9675 0.2625 1.3125 0.3375 ;
        RECT 0.8925 0.2625 0.9675 0.4875 ;
        RECT 0.6075 0.4125 0.8925 0.4875 ;
        VIA 0.9300 0.3525 VIA12_square ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 2.2800 0.3300 2.3850 0.4875 ;
        RECT 2.1900 0.4125 2.2800 0.4875 ;
        RECT 2.1150 0.4125 2.1900 0.6375 ;
        RECT 1.6500 0.5625 2.1150 0.6375 ;
        VIA 2.3325 0.4050 VIA12_square ;
        END
    END I1
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 3.8775 0.2175 3.9525 0.8325 ;
        RECT 3.8475 0.2175 3.8775 0.3825 ;
        RECT 3.8475 0.6675 3.8775 0.8325 ;
        END
    END Z
    PIN I0
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.2750 0.4350 1.3800 0.6375 ;
        RECT 0.8175 0.5625 1.2750 0.6375 ;
        VIA 1.3275 0.5100 VIA12_square ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 3.7350 -0.0750 3.9900 0.0750 ;
        RECT 3.6150 -0.0750 3.7350 0.2175 ;
        RECT 2.4675 -0.0750 3.6150 0.0750 ;
        RECT 2.3625 -0.0750 2.4675 0.2400 ;
        RECT 1.3950 -0.0750 2.3625 0.0750 ;
        RECT 1.2900 -0.0750 1.3950 0.2250 ;
        RECT 1.0050 -0.0750 1.2900 0.0750 ;
        RECT 0.8850 -0.0750 1.0050 0.2175 ;
        RECT 0.1425 -0.0750 0.8850 0.0750 ;
        RECT 0.0675 -0.0750 0.1425 0.2475 ;
        RECT 0.0000 -0.0750 0.0675 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 3.7200 0.9750 3.9900 1.1250 ;
        RECT 3.6450 0.7275 3.7200 1.1250 ;
        RECT 2.4750 0.9750 3.6450 1.1250 ;
        RECT 2.3550 0.8700 2.4750 1.1250 ;
        RECT 1.4400 0.9750 2.3550 1.1250 ;
        RECT 1.3350 0.8325 1.4400 1.1250 ;
        RECT 0.9750 0.9750 1.3350 1.1250 ;
        RECT 0.8700 0.8025 0.9750 1.1250 ;
        RECT 0.1425 0.9750 0.8700 1.1250 ;
        RECT 0.0675 0.7875 0.1425 1.1250 ;
        RECT 0.0000 0.9750 0.0675 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 3.8550 0.2700 3.9150 0.3300 ;
        RECT 3.8550 0.7200 3.9150 0.7800 ;
        RECT 3.7425 0.4875 3.8025 0.5475 ;
        RECT 3.6450 0.1575 3.7050 0.2175 ;
        RECT 3.6450 0.7575 3.7050 0.8175 ;
        RECT 3.2250 0.1725 3.2850 0.2325 ;
        RECT 3.2250 0.6750 3.2850 0.7350 ;
        RECT 3.1125 0.4800 3.1725 0.5400 ;
        RECT 3.0150 0.2100 3.0750 0.2700 ;
        RECT 3.0150 0.8100 3.0750 0.8700 ;
        RECT 2.9025 0.4050 2.9625 0.4650 ;
        RECT 2.8050 0.1875 2.8650 0.2475 ;
        RECT 2.8050 0.7650 2.8650 0.8250 ;
        RECT 2.5950 0.1800 2.6550 0.2400 ;
        RECT 2.5950 0.7875 2.6550 0.8475 ;
        RECT 2.4900 0.5625 2.5500 0.6225 ;
        RECT 2.3850 0.1575 2.4450 0.2175 ;
        RECT 2.3850 0.8700 2.4450 0.9300 ;
        RECT 2.2800 0.4800 2.3400 0.5400 ;
        RECT 2.0700 0.3300 2.1300 0.3900 ;
        RECT 2.0625 0.5700 2.1225 0.6300 ;
        RECT 1.9650 0.1575 2.0250 0.2175 ;
        RECT 1.9650 0.8325 2.0250 0.8925 ;
        RECT 1.8600 0.4875 1.9200 0.5475 ;
        RECT 1.7550 0.1575 1.8150 0.2175 ;
        RECT 1.7550 0.8325 1.8150 0.8925 ;
        RECT 1.6500 0.6300 1.7100 0.6900 ;
        RECT 1.5450 0.1575 1.6050 0.2175 ;
        RECT 1.4400 0.4800 1.5000 0.5400 ;
        RECT 1.3350 0.1350 1.3950 0.1950 ;
        RECT 1.3350 0.8700 1.3950 0.9300 ;
        RECT 1.2300 0.6450 1.2900 0.7050 ;
        RECT 1.1250 0.2775 1.1850 0.3375 ;
        RECT 1.1250 0.8325 1.1850 0.8925 ;
        RECT 0.9150 0.1575 0.9750 0.2175 ;
        RECT 0.9150 0.8325 0.9750 0.8925 ;
        RECT 0.8100 0.3300 0.8700 0.3900 ;
        RECT 0.6000 0.4125 0.6600 0.4725 ;
        RECT 0.6000 0.6525 0.6600 0.7125 ;
        RECT 0.4950 0.1575 0.5550 0.2175 ;
        RECT 0.4950 0.8325 0.5550 0.8925 ;
        RECT 0.3900 0.6525 0.4500 0.7125 ;
        RECT 0.3825 0.3300 0.4425 0.3900 ;
        RECT 0.1800 0.5925 0.2400 0.6525 ;
        RECT 0.0750 0.1575 0.1350 0.2175 ;
        RECT 0.0750 0.8175 0.1350 0.8775 ;
        LAYER M1 ;
        RECT 3.5700 0.4575 3.8025 0.5775 ;
        RECT 3.5400 0.2925 3.6375 0.3675 ;
        RECT 3.4950 0.4425 3.5700 0.9000 ;
        RECT 3.4575 0.1500 3.5400 0.3675 ;
        RECT 3.3825 0.4425 3.4950 0.5175 ;
        RECT 3.0900 0.8250 3.4950 0.9000 ;
        RECT 3.2025 0.1500 3.4575 0.2550 ;
        RECT 3.3075 0.5925 3.4200 0.7500 ;
        RECT 3.3075 0.3300 3.3825 0.5175 ;
        RECT 3.1275 0.3300 3.3075 0.4050 ;
        RECT 3.1875 0.6300 3.3075 0.7500 ;
        RECT 3.1125 0.4800 3.2025 0.5550 ;
        RECT 3.0525 0.1800 3.1275 0.4050 ;
        RECT 3.0375 0.4800 3.1125 0.6750 ;
        RECT 3.0150 0.7800 3.0900 0.9000 ;
        RECT 3.0150 0.1800 3.0525 0.3000 ;
        RECT 2.7900 0.6000 3.0375 0.6750 ;
        RECT 2.8575 0.3750 2.9625 0.4950 ;
        RECT 2.7300 0.1500 2.9400 0.3000 ;
        RECT 2.7300 0.7500 2.9400 0.9000 ;
        RECT 2.6550 0.3750 2.8575 0.4575 ;
        RECT 2.7225 0.5625 2.7900 0.6750 ;
        RECT 2.5875 0.5625 2.7225 0.6375 ;
        RECT 2.5500 0.1500 2.6550 0.4575 ;
        RECT 2.5500 0.7125 2.6550 0.8850 ;
        RECT 2.4600 0.5325 2.5875 0.6375 ;
        RECT 2.3850 0.7125 2.5500 0.7950 ;
        RECT 2.3850 0.3300 2.4750 0.4500 ;
        RECT 2.2800 0.3300 2.3850 0.6150 ;
        RECT 2.2050 0.4800 2.2800 0.6150 ;
        RECT 1.9350 0.1500 2.2725 0.2550 ;
        RECT 1.7925 0.3300 2.1750 0.4050 ;
        RECT 2.0550 0.4800 2.1300 0.6600 ;
        RECT 1.6725 0.4800 2.0550 0.5550 ;
        RECT 1.9800 0.8250 2.0550 0.9000 ;
        RECT 1.8300 0.6300 1.9800 0.9000 ;
        RECT 1.7325 0.1500 1.8600 0.2550 ;
        RECT 1.7250 0.8250 1.8300 0.9000 ;
        RECT 1.5825 0.6300 1.7550 0.7500 ;
        RECT 1.5000 0.1500 1.7325 0.2250 ;
        RECT 1.5975 0.3000 1.6725 0.5550 ;
        RECT 1.2000 0.3000 1.5975 0.3750 ;
        RECT 1.3200 0.6525 1.5825 0.7500 ;
        RECT 1.3650 0.4500 1.5225 0.5775 ;
        RECT 1.2525 0.4500 1.3650 0.5700 ;
        RECT 1.2000 0.6450 1.3200 0.7500 ;
        RECT 1.1250 0.8250 1.2225 0.9000 ;
        RECT 1.1775 0.2100 1.2000 0.3750 ;
        RECT 1.1250 0.2100 1.1775 0.5700 ;
        RECT 1.1025 0.2100 1.1250 0.9000 ;
        RECT 1.0500 0.4875 1.1025 0.9000 ;
        RECT 0.6900 0.4875 1.0500 0.5775 ;
        RECT 0.7650 0.2925 1.0275 0.4125 ;
        RECT 0.7950 0.6525 0.9450 0.7275 ;
        RECT 0.7200 0.6525 0.7950 0.8325 ;
        RECT 0.5550 0.6525 0.7200 0.7425 ;
        RECT 0.5700 0.4125 0.6900 0.5775 ;
        RECT 0.5175 0.1500 0.6825 0.3375 ;
        RECT 0.2475 0.8175 0.6150 0.9000 ;
        RECT 0.4500 0.5025 0.5700 0.5775 ;
        RECT 0.4650 0.1500 0.5175 0.2250 ;
        RECT 0.3300 0.5025 0.4500 0.7425 ;
        RECT 0.3600 0.3000 0.4425 0.4275 ;
        RECT 0.2175 0.1500 0.3600 0.4275 ;
        LAYER VIA1 ;
        RECT 3.5025 0.2925 3.5775 0.3675 ;
        RECT 3.2325 0.6600 3.3075 0.7350 ;
        RECT 2.8125 0.8100 2.8875 0.8850 ;
        RECT 2.7975 0.2100 2.8725 0.2850 ;
        RECT 2.6325 0.3750 2.7075 0.4500 ;
        RECT 2.5350 0.7125 2.6100 0.7875 ;
        RECT 2.0100 0.1575 2.0850 0.2325 ;
        RECT 1.8675 0.7125 1.9425 0.7875 ;
        RECT 0.5625 0.2625 0.6375 0.3375 ;
        RECT 0.3975 0.8175 0.4725 0.8925 ;
        LAYER M2 ;
        RECT 3.5025 0.2925 3.6225 0.3675 ;
        RECT 3.4275 0.2925 3.5025 0.9375 ;
        RECT 2.9250 0.8625 3.4275 0.9375 ;
        RECT 3.1875 0.6450 3.3525 0.7500 ;
        RECT 2.8725 0.6450 3.1875 0.7200 ;
        RECT 2.7750 0.7950 2.9250 0.9375 ;
        RECT 2.7975 0.1650 2.8725 0.7200 ;
        RECT 2.5425 0.1650 2.7975 0.2400 ;
        RECT 0.4725 0.8625 2.7750 0.9375 ;
        RECT 2.7000 0.3375 2.7225 0.4875 ;
        RECT 2.6175 0.3375 2.7000 0.7875 ;
        RECT 2.4900 0.7125 2.6175 0.7875 ;
        RECT 2.4675 0.1125 2.5425 0.6375 ;
        RECT 2.1000 0.1125 2.4675 0.1875 ;
        RECT 2.3400 0.5625 2.4675 0.6375 ;
        RECT 2.2650 0.5625 2.3400 0.7875 ;
        RECT 1.8225 0.7125 2.2650 0.7875 ;
        RECT 1.9950 0.1125 2.1000 0.2775 ;
        RECT 0.4725 0.2625 0.6825 0.3375 ;
        RECT 0.3975 0.2625 0.4725 0.9375 ;
    END
END MUX4_1010


MACRO ND2_0001
    CLASS CORE ;
    FOREIGN ND2_0001 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.4700 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 0.6075 0.7125 1.1025 0.7875 ;
        RECT 0.5025 0.2700 0.6075 0.7875 ;
        VIA 0.5550 0.3525 VIA12_square ;
        VIA 0.5550 0.7050 VIA12_square ;
        END
    END ZN
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.3275 0.4125 1.4025 0.6825 ;
        RECT 0.7800 0.4125 1.3275 0.5250 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1575 0.4800 0.6900 0.5850 ;
        RECT 0.0525 0.3675 0.1575 0.6825 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.2150 -0.0750 1.4700 0.0750 ;
        RECT 1.0950 -0.0750 1.2150 0.1875 ;
        RECT 0.0000 -0.0750 1.0950 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.4175 0.9750 1.4700 1.1250 ;
        RECT 1.3125 0.7875 1.4175 1.1250 ;
        RECT 0.9975 0.9750 1.3125 1.1250 ;
        RECT 0.8925 0.8250 0.9975 1.1250 ;
        RECT 0.5775 0.9750 0.8925 1.1250 ;
        RECT 0.4725 0.8250 0.5775 1.1250 ;
        RECT 0.1575 0.9750 0.4725 1.1250 ;
        RECT 0.0525 0.7875 0.1575 1.1250 ;
        RECT 0.0000 0.9750 0.0525 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.3350 0.2100 1.3950 0.2700 ;
        RECT 1.3350 0.8175 1.3950 0.8775 ;
        RECT 1.2300 0.4650 1.2900 0.5250 ;
        RECT 1.1250 0.1275 1.1850 0.1875 ;
        RECT 1.1250 0.7725 1.1850 0.8325 ;
        RECT 1.0200 0.4650 1.0800 0.5250 ;
        RECT 0.9150 0.2700 0.9750 0.3300 ;
        RECT 0.9150 0.8550 0.9750 0.9150 ;
        RECT 0.8100 0.4650 0.8700 0.5250 ;
        RECT 0.7050 0.6750 0.7650 0.7350 ;
        RECT 0.6000 0.4800 0.6600 0.5400 ;
        RECT 0.4950 0.1575 0.5550 0.2175 ;
        RECT 0.4950 0.8550 0.5550 0.9150 ;
        RECT 0.3900 0.4800 0.4500 0.5400 ;
        RECT 0.2850 0.3000 0.3450 0.3600 ;
        RECT 0.2850 0.7800 0.3450 0.8400 ;
        RECT 0.1800 0.4800 0.2400 0.5400 ;
        RECT 0.0750 0.1800 0.1350 0.2400 ;
        RECT 0.0750 0.8175 0.1350 0.8775 ;
        LAYER M1 ;
        RECT 1.3275 0.1800 1.4025 0.3375 ;
        RECT 0.8100 0.2625 1.3275 0.3375 ;
        RECT 1.1175 0.6675 1.1925 0.8700 ;
        RECT 0.3525 0.6675 1.1175 0.7425 ;
        RECT 0.7350 0.1500 0.8100 0.3375 ;
        RECT 0.1575 0.1500 0.7350 0.2250 ;
        RECT 0.2550 0.3000 0.6525 0.4050 ;
        RECT 0.2775 0.6675 0.3525 0.8700 ;
        RECT 0.0525 0.1500 0.1575 0.2700 ;
    END
END ND2_0001


MACRO ND2_0010
    CLASS CORE ;
    FOREIGN ND2_0010 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.4100 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 1.5225 0.2925 1.6800 0.4125 ;
        RECT 1.5225 0.6450 1.6800 0.7650 ;
        RECT 1.2075 0.2925 1.5225 0.7650 ;
        RECT 1.0500 0.2925 1.2075 0.4125 ;
        RECT 1.0500 0.6450 1.2075 0.7650 ;
        VIA 1.5225 0.3525 VIA12_slot ;
        VIA 1.5225 0.7050 VIA12_slot ;
        VIA 1.2075 0.3525 VIA12_slot ;
        VIA 1.2075 0.7050 VIA12_slot ;
        END
    END ZN
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 4.0725 0.4125 4.2375 0.6375 ;
        RECT 1.8300 0.4125 4.0725 0.5250 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1575 0.4800 1.7400 0.5850 ;
        RECT 0.0525 0.3675 0.1575 0.6825 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 4.1550 -0.0750 4.4100 0.0750 ;
        RECT 4.0350 -0.0750 4.1550 0.1875 ;
        RECT 3.7350 -0.0750 4.0350 0.0750 ;
        RECT 3.6150 -0.0750 3.7350 0.1875 ;
        RECT 3.3150 -0.0750 3.6150 0.0750 ;
        RECT 3.1950 -0.0750 3.3150 0.1875 ;
        RECT 2.8950 -0.0750 3.1950 0.0750 ;
        RECT 2.7750 -0.0750 2.8950 0.1875 ;
        RECT 2.4750 -0.0750 2.7750 0.0750 ;
        RECT 2.3550 -0.0750 2.4750 0.1875 ;
        RECT 2.0550 -0.0750 2.3550 0.0750 ;
        RECT 1.9350 -0.0750 2.0550 0.1875 ;
        RECT 0.0000 -0.0750 1.9350 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 4.3425 0.9750 4.4100 1.1250 ;
        RECT 4.2675 0.7800 4.3425 1.1250 ;
        RECT 3.9450 0.9750 4.2675 1.1250 ;
        RECT 3.8250 0.8625 3.9450 1.1250 ;
        RECT 3.5250 0.9750 3.8250 1.1250 ;
        RECT 3.4050 0.8625 3.5250 1.1250 ;
        RECT 3.1050 0.9750 3.4050 1.1250 ;
        RECT 2.9850 0.8625 3.1050 1.1250 ;
        RECT 2.6850 0.9750 2.9850 1.1250 ;
        RECT 2.5650 0.8625 2.6850 1.1250 ;
        RECT 2.2650 0.9750 2.5650 1.1250 ;
        RECT 2.1450 0.8625 2.2650 1.1250 ;
        RECT 1.8450 0.9750 2.1450 1.1250 ;
        RECT 1.7250 0.8625 1.8450 1.1250 ;
        RECT 1.4250 0.9750 1.7250 1.1250 ;
        RECT 1.3050 0.8625 1.4250 1.1250 ;
        RECT 1.0050 0.9750 1.3050 1.1250 ;
        RECT 0.8850 0.8625 1.0050 1.1250 ;
        RECT 0.5850 0.9750 0.8850 1.1250 ;
        RECT 0.4650 0.8625 0.5850 1.1250 ;
        RECT 0.1575 0.9750 0.4650 1.1250 ;
        RECT 0.0525 0.7875 0.1575 1.1250 ;
        RECT 0.0000 0.9750 0.0525 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 4.2750 0.2100 4.3350 0.2700 ;
        RECT 4.2750 0.8325 4.3350 0.8925 ;
        RECT 4.1700 0.4650 4.2300 0.5250 ;
        RECT 4.0650 0.1275 4.1250 0.1875 ;
        RECT 4.0650 0.8175 4.1250 0.8775 ;
        RECT 3.9600 0.4650 4.0200 0.5250 ;
        RECT 3.8550 0.2700 3.9150 0.3300 ;
        RECT 3.8550 0.8625 3.9150 0.9225 ;
        RECT 3.7500 0.4650 3.8100 0.5250 ;
        RECT 3.6450 0.1275 3.7050 0.1875 ;
        RECT 3.6450 0.8175 3.7050 0.8775 ;
        RECT 3.5400 0.4650 3.6000 0.5250 ;
        RECT 3.4350 0.2700 3.4950 0.3300 ;
        RECT 3.4350 0.8625 3.4950 0.9225 ;
        RECT 3.3300 0.4650 3.3900 0.5250 ;
        RECT 3.2250 0.1275 3.2850 0.1875 ;
        RECT 3.2250 0.8175 3.2850 0.8775 ;
        RECT 3.1200 0.4650 3.1800 0.5250 ;
        RECT 3.0150 0.2700 3.0750 0.3300 ;
        RECT 3.0150 0.8625 3.0750 0.9225 ;
        RECT 2.9100 0.4650 2.9700 0.5250 ;
        RECT 2.8050 0.1275 2.8650 0.1875 ;
        RECT 2.8050 0.8175 2.8650 0.8775 ;
        RECT 2.7000 0.4650 2.7600 0.5250 ;
        RECT 2.5950 0.2700 2.6550 0.3300 ;
        RECT 2.5950 0.8625 2.6550 0.9225 ;
        RECT 2.4900 0.4650 2.5500 0.5250 ;
        RECT 2.3850 0.1275 2.4450 0.1875 ;
        RECT 2.3850 0.6975 2.4450 0.7575 ;
        RECT 2.2800 0.4650 2.3400 0.5250 ;
        RECT 2.1750 0.2700 2.2350 0.3300 ;
        RECT 2.1750 0.8625 2.2350 0.9225 ;
        RECT 2.0700 0.4650 2.1300 0.5250 ;
        RECT 1.9650 0.1275 2.0250 0.1875 ;
        RECT 1.9650 0.6975 2.0250 0.7575 ;
        RECT 1.8600 0.4650 1.9200 0.5250 ;
        RECT 1.7550 0.1575 1.8150 0.2175 ;
        RECT 1.7550 0.8625 1.8150 0.9225 ;
        RECT 1.6500 0.4800 1.7100 0.5400 ;
        RECT 1.5450 0.3000 1.6050 0.3600 ;
        RECT 1.5450 0.6975 1.6050 0.7575 ;
        RECT 1.4400 0.4800 1.5000 0.5400 ;
        RECT 1.3350 0.1575 1.3950 0.2175 ;
        RECT 1.3350 0.8625 1.3950 0.9225 ;
        RECT 1.2300 0.4800 1.2900 0.5400 ;
        RECT 1.1250 0.3000 1.1850 0.3600 ;
        RECT 1.1250 0.6975 1.1850 0.7575 ;
        RECT 1.0200 0.4800 1.0800 0.5400 ;
        RECT 0.9150 0.1575 0.9750 0.2175 ;
        RECT 0.9150 0.8625 0.9750 0.9225 ;
        RECT 0.2850 0.6975 0.3450 0.7575 ;
        RECT 0.1800 0.4800 0.2400 0.5400 ;
        RECT 0.0750 0.1800 0.1350 0.2400 ;
        RECT 0.0750 0.8175 0.1350 0.8775 ;
        RECT 0.8100 0.4800 0.8700 0.5400 ;
        RECT 0.7050 0.3000 0.7650 0.3600 ;
        RECT 0.7050 0.6975 0.7650 0.7575 ;
        RECT 0.6000 0.4800 0.6600 0.5400 ;
        RECT 0.4950 0.1575 0.5550 0.2175 ;
        RECT 0.4950 0.8625 0.5550 0.9225 ;
        RECT 0.3900 0.4800 0.4500 0.5400 ;
        RECT 0.2850 0.3000 0.3450 0.3600 ;
        LAYER M1 ;
        RECT 4.2675 0.1800 4.3425 0.3375 ;
        RECT 1.8525 0.2625 4.2675 0.3375 ;
        RECT 4.0425 0.7125 4.1475 0.9000 ;
        RECT 3.9975 0.7125 4.0425 0.7875 ;
        RECT 3.7275 0.6675 3.9975 0.7875 ;
        RECT 3.6225 0.6675 3.7275 0.9000 ;
        RECT 3.3075 0.6675 3.6225 0.7875 ;
        RECT 3.2025 0.6675 3.3075 0.9000 ;
        RECT 2.8875 0.6675 3.2025 0.7875 ;
        RECT 2.7825 0.6675 2.8875 0.9000 ;
        RECT 0.2775 0.6675 2.7825 0.7875 ;
        RECT 1.7775 0.1500 1.8525 0.3375 ;
        RECT 0.1575 0.1500 1.7775 0.2250 ;
        RECT 0.2550 0.3000 1.7025 0.4050 ;
        RECT 0.0525 0.1500 0.1575 0.2700 ;
        LAYER M2 ;
        RECT 1.5525 0.2925 1.6800 0.4125 ;
        RECT 1.5525 0.6450 1.6800 0.7650 ;
        RECT 1.0500 0.2925 1.1775 0.4125 ;
        RECT 1.0500 0.6450 1.1775 0.7650 ;
    END
END ND2_0010


MACRO ND2_0011
    CLASS CORE ;
    FOREIGN ND2_0011 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.0500 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.6975 0.7125 0.7725 0.8325 ;
        RECT 0.2925 0.7125 0.6975 0.7875 ;
        RECT 0.2550 0.3000 0.3675 0.4050 ;
        RECT 0.2325 0.6750 0.2925 0.7875 ;
        RECT 0.1125 0.3300 0.2550 0.4050 ;
        RECT 0.1125 0.6750 0.2325 0.7575 ;
        RECT 0.0375 0.3300 0.1125 0.7575 ;
        END
    END ZN
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.9075 0.4125 1.0125 0.6825 ;
        RECT 0.6075 0.4125 0.9075 0.5625 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.4575 0.3675 0.5325 0.6375 ;
        RECT 0.3675 0.4800 0.4575 0.6375 ;
        RECT 0.1875 0.4800 0.3675 0.6000 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.7950 -0.0750 1.0500 0.0750 ;
        RECT 0.6750 -0.0750 0.7950 0.1875 ;
        RECT 0.0000 -0.0750 0.6750 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.9825 0.9750 1.0500 1.1250 ;
        RECT 0.9075 0.8025 0.9825 1.1250 ;
        RECT 0.5850 0.9750 0.9075 1.1250 ;
        RECT 0.4650 0.8625 0.5850 1.1250 ;
        RECT 0.1650 0.9750 0.4650 1.1250 ;
        RECT 0.0450 0.8325 0.1650 1.1250 ;
        RECT 0.0000 0.9750 0.0450 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 0.9150 0.2100 0.9750 0.2700 ;
        RECT 0.9150 0.8325 0.9750 0.8925 ;
        RECT 0.8100 0.4650 0.8700 0.5250 ;
        RECT 0.7050 0.1200 0.7650 0.1800 ;
        RECT 0.7050 0.7425 0.7650 0.8025 ;
        RECT 0.6075 0.4650 0.6675 0.5250 ;
        RECT 0.4950 0.1725 0.5550 0.2325 ;
        RECT 0.4950 0.8700 0.5550 0.9300 ;
        RECT 0.3900 0.5100 0.4500 0.5700 ;
        RECT 0.2850 0.3225 0.3450 0.3825 ;
        RECT 0.2850 0.7200 0.3450 0.7800 ;
        RECT 0.1875 0.5100 0.2475 0.5700 ;
        RECT 0.0750 0.1725 0.1350 0.2325 ;
        RECT 0.0750 0.8325 0.1350 0.8925 ;
        LAYER M1 ;
        RECT 0.8925 0.1800 0.9975 0.3375 ;
        RECT 0.6900 0.2625 0.8925 0.3375 ;
        RECT 0.4350 0.1500 0.5850 0.2550 ;
        RECT 0.1650 0.1500 0.4350 0.2250 ;
        RECT 0.0450 0.1500 0.1650 0.2550 ;
        LAYER VIA1 ;
        RECT 0.7350 0.2625 0.8100 0.3375 ;
        RECT 0.4725 0.1650 0.5475 0.2400 ;
        LAYER M2 ;
        RECT 0.7200 0.2625 0.8850 0.3375 ;
        RECT 0.6450 0.1650 0.7200 0.3375 ;
        RECT 0.3975 0.1650 0.6450 0.2400 ;
    END
END ND2_0011


MACRO ND2_0100
    CLASS CORE ;
    FOREIGN ND2_0100 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.5700 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 1.1025 0.2925 1.2600 0.4125 ;
        RECT 1.1025 0.6450 1.2600 0.7650 ;
        RECT 0.7875 0.2925 1.1025 0.7650 ;
        RECT 0.6300 0.2925 0.7875 0.4125 ;
        RECT 0.6300 0.6450 0.7875 0.7650 ;
        VIA 1.1025 0.3525 VIA12_slot ;
        VIA 1.1025 0.7050 VIA12_slot ;
        VIA 0.7875 0.3525 VIA12_slot ;
        VIA 0.7875 0.7050 VIA12_slot ;
        END
    END ZN
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 3.4275 0.4125 3.5025 0.6825 ;
        RECT 1.8300 0.4125 3.4275 0.5250 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1575 0.4800 1.7400 0.5850 ;
        RECT 0.0525 0.3675 0.1575 0.6825 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 3.3150 -0.0750 3.5700 0.0750 ;
        RECT 3.1950 -0.0750 3.3150 0.1875 ;
        RECT 2.8950 -0.0750 3.1950 0.0750 ;
        RECT 2.7750 -0.0750 2.8950 0.1875 ;
        RECT 2.4750 -0.0750 2.7750 0.0750 ;
        RECT 2.3550 -0.0750 2.4750 0.1875 ;
        RECT 2.0550 -0.0750 2.3550 0.0750 ;
        RECT 1.9350 -0.0750 2.0550 0.1875 ;
        RECT 0.0000 -0.0750 1.9350 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 3.5175 0.9750 3.5700 1.1250 ;
        RECT 3.4125 0.7875 3.5175 1.1250 ;
        RECT 3.0975 0.9750 3.4125 1.1250 ;
        RECT 2.9925 0.8250 3.0975 1.1250 ;
        RECT 2.6775 0.9750 2.9925 1.1250 ;
        RECT 2.5725 0.8250 2.6775 1.1250 ;
        RECT 2.2575 0.9750 2.5725 1.1250 ;
        RECT 2.1525 0.8250 2.2575 1.1250 ;
        RECT 1.8375 0.9750 2.1525 1.1250 ;
        RECT 1.7325 0.8250 1.8375 1.1250 ;
        RECT 1.4175 0.9750 1.7325 1.1250 ;
        RECT 1.3125 0.8250 1.4175 1.1250 ;
        RECT 0.9975 0.9750 1.3125 1.1250 ;
        RECT 0.8925 0.8250 0.9975 1.1250 ;
        RECT 0.5775 0.9750 0.8925 1.1250 ;
        RECT 0.4725 0.8250 0.5775 1.1250 ;
        RECT 0.1575 0.9750 0.4725 1.1250 ;
        RECT 0.0525 0.7875 0.1575 1.1250 ;
        RECT 0.0000 0.9750 0.0525 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 3.4350 0.2100 3.4950 0.2700 ;
        RECT 3.4350 0.8175 3.4950 0.8775 ;
        RECT 3.3300 0.4650 3.3900 0.5250 ;
        RECT 3.2250 0.1275 3.2850 0.1875 ;
        RECT 3.2250 0.7725 3.2850 0.8325 ;
        RECT 3.1200 0.4650 3.1800 0.5250 ;
        RECT 3.0150 0.2700 3.0750 0.3300 ;
        RECT 3.0150 0.8550 3.0750 0.9150 ;
        RECT 2.9100 0.4650 2.9700 0.5250 ;
        RECT 2.8050 0.1275 2.8650 0.1875 ;
        RECT 2.8050 0.6750 2.8650 0.7350 ;
        RECT 2.7000 0.4650 2.7600 0.5250 ;
        RECT 2.5950 0.2700 2.6550 0.3300 ;
        RECT 2.5950 0.8550 2.6550 0.9150 ;
        RECT 2.4900 0.4650 2.5500 0.5250 ;
        RECT 2.3850 0.1275 2.4450 0.1875 ;
        RECT 2.3850 0.6750 2.4450 0.7350 ;
        RECT 2.2800 0.4650 2.3400 0.5250 ;
        RECT 2.1750 0.2700 2.2350 0.3300 ;
        RECT 2.1750 0.8550 2.2350 0.9150 ;
        RECT 2.0700 0.4650 2.1300 0.5250 ;
        RECT 1.9650 0.1275 2.0250 0.1875 ;
        RECT 1.9650 0.6750 2.0250 0.7350 ;
        RECT 1.8600 0.4650 1.9200 0.5250 ;
        RECT 1.7550 0.1575 1.8150 0.2175 ;
        RECT 1.7550 0.8550 1.8150 0.9150 ;
        RECT 1.6500 0.4800 1.7100 0.5400 ;
        RECT 1.5450 0.3000 1.6050 0.3600 ;
        RECT 0.9150 0.1575 0.9750 0.2175 ;
        RECT 0.9150 0.8550 0.9750 0.9150 ;
        RECT 0.8100 0.4800 0.8700 0.5400 ;
        RECT 0.7050 0.3000 0.7650 0.3600 ;
        RECT 0.7050 0.6750 0.7650 0.7350 ;
        RECT 0.6000 0.4800 0.6600 0.5400 ;
        RECT 0.4950 0.1575 0.5550 0.2175 ;
        RECT 0.4950 0.8550 0.5550 0.9150 ;
        RECT 0.3900 0.4800 0.4500 0.5400 ;
        RECT 0.2850 0.3000 0.3450 0.3600 ;
        RECT 0.2850 0.7800 0.3450 0.8400 ;
        RECT 0.1800 0.4800 0.2400 0.5400 ;
        RECT 0.0750 0.1800 0.1350 0.2400 ;
        RECT 0.0750 0.8175 0.1350 0.8775 ;
        RECT 1.5450 0.6750 1.6050 0.7350 ;
        RECT 1.4400 0.4800 1.5000 0.5400 ;
        RECT 1.3350 0.1575 1.3950 0.2175 ;
        RECT 1.3350 0.8550 1.3950 0.9150 ;
        RECT 1.2300 0.4800 1.2900 0.5400 ;
        RECT 1.1250 0.3000 1.1850 0.3600 ;
        RECT 1.1250 0.6750 1.1850 0.7350 ;
        RECT 1.0200 0.4800 1.0800 0.5400 ;
        LAYER M1 ;
        RECT 3.4275 0.1800 3.5025 0.3375 ;
        RECT 1.8525 0.2625 3.4275 0.3375 ;
        RECT 3.2175 0.6675 3.2925 0.8700 ;
        RECT 0.3525 0.6675 3.2175 0.7425 ;
        RECT 1.7775 0.1500 1.8525 0.3375 ;
        RECT 0.1575 0.1500 1.7775 0.2250 ;
        RECT 0.2550 0.3000 1.7025 0.4050 ;
        RECT 0.2775 0.6675 0.3525 0.8700 ;
        RECT 0.0525 0.1500 0.1575 0.2700 ;
        LAYER M2 ;
        RECT 1.1325 0.2925 1.2600 0.4125 ;
        RECT 1.1325 0.6450 1.2600 0.7650 ;
        RECT 0.6300 0.2925 0.7575 0.4125 ;
        RECT 0.6300 0.6450 0.7575 0.7650 ;
    END
END ND2_0100


MACRO ND2_0101
    CLASS CORE ;
    FOREIGN ND2_0101 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.2500 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 1.9425 0.2925 2.1000 0.4125 ;
        RECT 1.9425 0.6450 2.1000 0.7650 ;
        RECT 1.6275 0.2925 1.9425 0.7650 ;
        RECT 1.4700 0.2925 1.6275 0.4125 ;
        RECT 1.4700 0.6450 1.6275 0.7650 ;
        VIA 1.9425 0.3525 VIA12_slot ;
        VIA 1.9425 0.7050 VIA12_slot ;
        VIA 1.6275 0.3525 VIA12_slot ;
        VIA 1.6275 0.7050 VIA12_slot ;
        END
    END ZN
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 5.1075 0.4125 5.1825 0.6825 ;
        RECT 2.6700 0.4125 5.1075 0.5250 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1575 0.4800 2.5800 0.5850 ;
        RECT 0.0525 0.3675 0.1575 0.6825 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 4.9950 -0.0750 5.2500 0.0750 ;
        RECT 4.8750 -0.0750 4.9950 0.1875 ;
        RECT 4.5750 -0.0750 4.8750 0.0750 ;
        RECT 4.4550 -0.0750 4.5750 0.1875 ;
        RECT 4.1550 -0.0750 4.4550 0.0750 ;
        RECT 4.0350 -0.0750 4.1550 0.1875 ;
        RECT 3.7350 -0.0750 4.0350 0.0750 ;
        RECT 3.6150 -0.0750 3.7350 0.1875 ;
        RECT 3.3150 -0.0750 3.6150 0.0750 ;
        RECT 3.1950 -0.0750 3.3150 0.1875 ;
        RECT 2.8950 -0.0750 3.1950 0.0750 ;
        RECT 2.7750 -0.0750 2.8950 0.1875 ;
        RECT 0.0000 -0.0750 2.7750 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 5.1975 0.9750 5.2500 1.1250 ;
        RECT 5.0925 0.7875 5.1975 1.1250 ;
        RECT 4.7775 0.9750 5.0925 1.1250 ;
        RECT 4.6725 0.8250 4.7775 1.1250 ;
        RECT 4.3575 0.9750 4.6725 1.1250 ;
        RECT 4.2525 0.8250 4.3575 1.1250 ;
        RECT 3.9375 0.9750 4.2525 1.1250 ;
        RECT 3.8325 0.8250 3.9375 1.1250 ;
        RECT 3.5175 0.9750 3.8325 1.1250 ;
        RECT 3.4125 0.8250 3.5175 1.1250 ;
        RECT 3.0975 0.9750 3.4125 1.1250 ;
        RECT 2.9925 0.8250 3.0975 1.1250 ;
        RECT 2.6775 0.9750 2.9925 1.1250 ;
        RECT 2.5725 0.8250 2.6775 1.1250 ;
        RECT 2.2575 0.9750 2.5725 1.1250 ;
        RECT 2.1525 0.8250 2.2575 1.1250 ;
        RECT 1.8375 0.9750 2.1525 1.1250 ;
        RECT 1.7325 0.8250 1.8375 1.1250 ;
        RECT 1.4175 0.9750 1.7325 1.1250 ;
        RECT 1.3125 0.8250 1.4175 1.1250 ;
        RECT 0.9975 0.9750 1.3125 1.1250 ;
        RECT 0.8925 0.8325 0.9975 1.1250 ;
        RECT 0.5775 0.9750 0.8925 1.1250 ;
        RECT 0.4725 0.8250 0.5775 1.1250 ;
        RECT 0.1575 0.9750 0.4725 1.1250 ;
        RECT 0.0525 0.7875 0.1575 1.1250 ;
        RECT 0.0000 0.9750 0.0525 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 5.1150 0.2100 5.1750 0.2700 ;
        RECT 5.1150 0.8175 5.1750 0.8775 ;
        RECT 5.0100 0.4650 5.0700 0.5250 ;
        RECT 4.9050 0.1275 4.9650 0.1875 ;
        RECT 4.9050 0.7725 4.9650 0.8325 ;
        RECT 4.8000 0.4650 4.8600 0.5250 ;
        RECT 4.6950 0.2700 4.7550 0.3300 ;
        RECT 4.6950 0.8550 4.7550 0.9150 ;
        RECT 4.5900 0.4650 4.6500 0.5250 ;
        RECT 4.4850 0.1275 4.5450 0.1875 ;
        RECT 4.4850 0.6750 4.5450 0.7350 ;
        RECT 4.3800 0.4650 4.4400 0.5250 ;
        RECT 4.2750 0.2700 4.3350 0.3300 ;
        RECT 4.2750 0.8550 4.3350 0.9150 ;
        RECT 4.1700 0.4650 4.2300 0.5250 ;
        RECT 4.0650 0.1275 4.1250 0.1875 ;
        RECT 4.0650 0.6750 4.1250 0.7350 ;
        RECT 3.9600 0.4650 4.0200 0.5250 ;
        RECT 3.8550 0.2700 3.9150 0.3300 ;
        RECT 3.8550 0.8550 3.9150 0.9150 ;
        RECT 3.7500 0.4650 3.8100 0.5250 ;
        RECT 3.6450 0.1275 3.7050 0.1875 ;
        RECT 3.6450 0.6750 3.7050 0.7350 ;
        RECT 3.5400 0.4650 3.6000 0.5250 ;
        RECT 3.4350 0.2700 3.4950 0.3300 ;
        RECT 3.4350 0.8550 3.4950 0.9150 ;
        RECT 3.3300 0.4650 3.3900 0.5250 ;
        RECT 3.2250 0.1275 3.2850 0.1875 ;
        RECT 3.2250 0.6750 3.2850 0.7350 ;
        RECT 3.1200 0.4650 3.1800 0.5250 ;
        RECT 3.0150 0.2700 3.0750 0.3300 ;
        RECT 3.0150 0.8550 3.0750 0.9150 ;
        RECT 2.9100 0.4650 2.9700 0.5250 ;
        RECT 2.8050 0.1275 2.8650 0.1875 ;
        RECT 2.8050 0.6750 2.8650 0.7350 ;
        RECT 2.7000 0.4650 2.7600 0.5250 ;
        RECT 2.5950 0.1575 2.6550 0.2175 ;
        RECT 2.5950 0.8550 2.6550 0.9150 ;
        RECT 2.4900 0.4800 2.5500 0.5400 ;
        RECT 2.3850 0.3000 2.4450 0.3600 ;
        RECT 2.3850 0.6750 2.4450 0.7350 ;
        RECT 2.2800 0.4800 2.3400 0.5400 ;
        RECT 2.1750 0.1575 2.2350 0.2175 ;
        RECT 2.1750 0.8550 2.2350 0.9150 ;
        RECT 2.0700 0.4800 2.1300 0.5400 ;
        RECT 1.9650 0.3000 2.0250 0.3600 ;
        RECT 1.9650 0.6750 2.0250 0.7350 ;
        RECT 1.8600 0.4800 1.9200 0.5400 ;
        RECT 1.7550 0.1575 1.8150 0.2175 ;
        RECT 1.7550 0.8550 1.8150 0.9150 ;
        RECT 1.6500 0.4800 1.7100 0.5400 ;
        RECT 1.5450 0.3000 1.6050 0.3600 ;
        RECT 1.5450 0.6750 1.6050 0.7350 ;
        RECT 1.4400 0.4800 1.5000 0.5400 ;
        RECT 1.3350 0.1575 1.3950 0.2175 ;
        RECT 1.3350 0.8550 1.3950 0.9150 ;
        RECT 1.2300 0.4800 1.2900 0.5400 ;
        RECT 1.1250 0.3000 1.1850 0.3600 ;
        RECT 0.4950 0.1575 0.5550 0.2175 ;
        RECT 0.4950 0.8550 0.5550 0.9150 ;
        RECT 0.3900 0.4800 0.4500 0.5400 ;
        RECT 0.2850 0.3000 0.3450 0.3600 ;
        RECT 0.2850 0.7800 0.3450 0.8400 ;
        RECT 0.1800 0.4800 0.2400 0.5400 ;
        RECT 0.0750 0.1800 0.1350 0.2400 ;
        RECT 0.0750 0.8175 0.1350 0.8775 ;
        RECT 1.1250 0.6825 1.1850 0.7425 ;
        RECT 1.0200 0.4800 1.0800 0.5400 ;
        RECT 0.9150 0.1575 0.9750 0.2175 ;
        RECT 0.9150 0.8550 0.9750 0.9150 ;
        RECT 0.8100 0.4800 0.8700 0.5400 ;
        RECT 0.7050 0.3000 0.7650 0.3600 ;
        RECT 0.7050 0.6750 0.7650 0.7350 ;
        RECT 0.6000 0.4800 0.6600 0.5400 ;
        LAYER M1 ;
        RECT 5.1075 0.1800 5.1825 0.3375 ;
        RECT 2.6925 0.2625 5.1075 0.3375 ;
        RECT 4.8975 0.6675 4.9725 0.8700 ;
        RECT 0.3525 0.6675 4.8975 0.7425 ;
        RECT 2.6175 0.1500 2.6925 0.3375 ;
        RECT 0.1575 0.1500 2.6175 0.2250 ;
        RECT 0.2550 0.3000 2.5425 0.4050 ;
        RECT 0.2775 0.6675 0.3525 0.8700 ;
        RECT 0.0525 0.1500 0.1575 0.2700 ;
        LAYER M2 ;
        RECT 1.9725 0.2925 2.1000 0.4125 ;
        RECT 1.9725 0.6450 2.1000 0.7650 ;
        RECT 1.4700 0.2925 1.5975 0.4125 ;
        RECT 1.4700 0.6450 1.5975 0.7650 ;
    END
END ND2_0101


MACRO ND2_0111
    CLASS CORE ;
    FOREIGN ND2_0111 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.8900 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 0.3675 0.2925 0.6825 0.7650 ;
        VIA 0.5250 0.3525 VIA12_slot ;
        VIA 0.5250 0.7050 VIA12_slot ;
        END
    END ZN
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.7475 0.4125 1.8225 0.6825 ;
        RECT 0.9975 0.4125 1.7475 0.5250 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1575 0.4800 0.9000 0.5850 ;
        RECT 0.0525 0.3675 0.1575 0.6825 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.6350 -0.0750 1.8900 0.0750 ;
        RECT 1.5150 -0.0750 1.6350 0.1875 ;
        RECT 1.2150 -0.0750 1.5150 0.0750 ;
        RECT 1.0950 -0.0750 1.2150 0.1875 ;
        RECT 0.0000 -0.0750 1.0950 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.8375 0.9750 1.8900 1.1250 ;
        RECT 1.7325 0.7875 1.8375 1.1250 ;
        RECT 1.4175 0.9750 1.7325 1.1250 ;
        RECT 1.3125 0.8250 1.4175 1.1250 ;
        RECT 0.9975 0.9750 1.3125 1.1250 ;
        RECT 0.8925 0.8250 0.9975 1.1250 ;
        RECT 0.5775 0.9750 0.8925 1.1250 ;
        RECT 0.4725 0.8250 0.5775 1.1250 ;
        RECT 0.1575 0.9750 0.4725 1.1250 ;
        RECT 0.0525 0.7875 0.1575 1.1250 ;
        RECT 0.0000 0.9750 0.0525 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.7550 0.2100 1.8150 0.2700 ;
        RECT 1.7550 0.8175 1.8150 0.8775 ;
        RECT 1.6500 0.4650 1.7100 0.5250 ;
        RECT 1.5450 0.1275 1.6050 0.1875 ;
        RECT 1.5450 0.7725 1.6050 0.8325 ;
        RECT 1.4400 0.4650 1.5000 0.5250 ;
        RECT 1.3350 0.2700 1.3950 0.3300 ;
        RECT 1.3350 0.8550 1.3950 0.9150 ;
        RECT 1.2300 0.4650 1.2900 0.5250 ;
        RECT 1.1250 0.1275 1.1850 0.1875 ;
        RECT 1.1250 0.6750 1.1850 0.7350 ;
        RECT 1.0275 0.4650 1.0875 0.5250 ;
        RECT 0.9150 0.1575 0.9750 0.2175 ;
        RECT 0.9150 0.8550 0.9750 0.9150 ;
        RECT 0.8100 0.4800 0.8700 0.5400 ;
        RECT 0.7050 0.3000 0.7650 0.3600 ;
        RECT 0.7050 0.6750 0.7650 0.7350 ;
        RECT 0.6000 0.4800 0.6600 0.5400 ;
        RECT 0.4950 0.1575 0.5550 0.2175 ;
        RECT 0.4950 0.8550 0.5550 0.9150 ;
        RECT 0.3900 0.4800 0.4500 0.5400 ;
        RECT 0.2850 0.3000 0.3450 0.3600 ;
        RECT 0.2850 0.7800 0.3450 0.8400 ;
        RECT 0.1800 0.4800 0.2400 0.5400 ;
        RECT 0.0750 0.1800 0.1350 0.2400 ;
        RECT 0.0750 0.8175 0.1350 0.8775 ;
        LAYER M1 ;
        RECT 1.7475 0.1800 1.8225 0.3375 ;
        RECT 1.0200 0.2625 1.7475 0.3375 ;
        RECT 1.5375 0.6675 1.6125 0.8700 ;
        RECT 0.3525 0.6675 1.5375 0.7425 ;
        RECT 0.9450 0.1500 1.0200 0.3375 ;
        RECT 0.1575 0.1500 0.9450 0.2250 ;
        RECT 0.2550 0.3000 0.8625 0.4050 ;
        RECT 0.2775 0.6675 0.3525 0.8700 ;
        RECT 0.0525 0.1500 0.1575 0.2700 ;
    END
END ND2_0111


MACRO ND2_1000
    CLASS CORE ;
    FOREIGN ND2_1000 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.6300 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.5175 0.1500 0.5925 0.7425 ;
        RECT 0.4725 0.1500 0.5175 0.3675 ;
        RECT 0.3675 0.6675 0.5175 0.7425 ;
        RECT 0.2625 0.6675 0.3675 0.8925 ;
        END
    END ZN
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1425 0.4575 0.2325 0.5925 ;
        RECT 0.0675 0.3675 0.1425 0.6825 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.0825 0.2625 0.5475 0.3375 ;
        VIA 0.3300 0.3000 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.1425 -0.0750 0.6300 0.0750 ;
        RECT 0.0675 -0.0750 0.1425 0.2475 ;
        RECT 0.0000 -0.0750 0.0675 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.5925 0.9750 0.6300 1.1250 ;
        RECT 0.4575 0.8175 0.5925 1.1250 ;
        RECT 0.1425 0.9750 0.4575 1.1250 ;
        RECT 0.0675 0.8025 0.1425 1.1250 ;
        RECT 0.0000 0.9750 0.0675 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 0.4950 0.1725 0.5550 0.2325 ;
        RECT 0.4950 0.8325 0.5550 0.8925 ;
        RECT 0.3825 0.4875 0.4425 0.5475 ;
        RECT 0.2850 0.8100 0.3450 0.8700 ;
        RECT 0.1725 0.4875 0.2325 0.5475 ;
        RECT 0.0750 0.1575 0.1350 0.2175 ;
        RECT 0.0750 0.8325 0.1350 0.8925 ;
        LAYER M1 ;
        RECT 0.3825 0.4425 0.4425 0.5925 ;
        RECT 0.3075 0.2175 0.3825 0.5925 ;
        RECT 0.2775 0.2175 0.3075 0.3825 ;
    END
END ND2_1000


MACRO ND2_1010
    CLASS CORE ;
    FOREIGN ND2_1010 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.6300 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.5175 0.2175 0.5925 0.7425 ;
        RECT 0.4875 0.2175 0.5175 0.3825 ;
        RECT 0.3525 0.6675 0.5175 0.7425 ;
        RECT 0.2775 0.6675 0.3525 0.8325 ;
        END
    END ZN
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1425 0.4575 0.2325 0.5925 ;
        RECT 0.0675 0.3675 0.1425 0.6825 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.3825 0.4425 0.4425 0.5925 ;
        RECT 0.3075 0.2175 0.3825 0.5925 ;
        RECT 0.2775 0.2175 0.3075 0.3825 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.1425 -0.0750 0.6300 0.0750 ;
        RECT 0.0675 -0.0750 0.1425 0.2475 ;
        RECT 0.0000 -0.0750 0.0675 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.5925 0.9750 0.6300 1.1250 ;
        RECT 0.4575 0.8175 0.5925 1.1250 ;
        RECT 0.1425 0.9750 0.4575 1.1250 ;
        RECT 0.0675 0.8025 0.1425 1.1250 ;
        RECT 0.0000 0.9750 0.0675 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 0.4950 0.2700 0.5550 0.3300 ;
        RECT 0.4950 0.8325 0.5550 0.8925 ;
        RECT 0.3825 0.4875 0.4425 0.5475 ;
        RECT 0.2850 0.7275 0.3450 0.7875 ;
        RECT 0.1725 0.4875 0.2325 0.5475 ;
        RECT 0.0750 0.1575 0.1350 0.2175 ;
        RECT 0.0750 0.8325 0.1350 0.8925 ;
    END
END ND2_1010


MACRO ND2_1100
    CLASS CORE ;
    FOREIGN ND2_1100 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.9300 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 2.7825 0.2925 2.9400 0.4125 ;
        RECT 2.7825 0.6450 2.9400 0.7650 ;
        RECT 2.4675 0.2925 2.7825 0.7650 ;
        RECT 2.3100 0.2925 2.4675 0.4125 ;
        RECT 2.3100 0.6450 2.4675 0.7650 ;
        VIA 2.7825 0.3525 VIA12_slot ;
        VIA 2.7825 0.7050 VIA12_slot ;
        VIA 2.4675 0.3525 VIA12_slot ;
        VIA 2.4675 0.7050 VIA12_slot ;
        END
    END ZN
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 6.7875 0.4125 6.8625 0.6825 ;
        RECT 3.5100 0.4125 6.7875 0.5250 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1575 0.4800 3.4200 0.5850 ;
        RECT 0.0525 0.3675 0.1575 0.6825 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 6.6750 -0.0750 6.9300 0.0750 ;
        RECT 6.5550 -0.0750 6.6750 0.1875 ;
        RECT 6.2550 -0.0750 6.5550 0.0750 ;
        RECT 6.1350 -0.0750 6.2550 0.1875 ;
        RECT 5.8350 -0.0750 6.1350 0.0750 ;
        RECT 5.7150 -0.0750 5.8350 0.1875 ;
        RECT 5.4150 -0.0750 5.7150 0.0750 ;
        RECT 5.2950 -0.0750 5.4150 0.1875 ;
        RECT 4.9950 -0.0750 5.2950 0.0750 ;
        RECT 4.8750 -0.0750 4.9950 0.1875 ;
        RECT 4.5750 -0.0750 4.8750 0.0750 ;
        RECT 4.4550 -0.0750 4.5750 0.1875 ;
        RECT 4.1550 -0.0750 4.4550 0.0750 ;
        RECT 4.0350 -0.0750 4.1550 0.1875 ;
        RECT 3.7350 -0.0750 4.0350 0.0750 ;
        RECT 3.6150 -0.0750 3.7350 0.1875 ;
        RECT 0.0000 -0.0750 3.6150 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 6.8775 0.9750 6.9300 1.1250 ;
        RECT 6.7725 0.7875 6.8775 1.1250 ;
        RECT 6.4575 0.9750 6.7725 1.1250 ;
        RECT 6.3525 0.8250 6.4575 1.1250 ;
        RECT 6.0375 0.9750 6.3525 1.1250 ;
        RECT 5.9325 0.8325 6.0375 1.1250 ;
        RECT 5.6175 0.9750 5.9325 1.1250 ;
        RECT 5.5125 0.8250 5.6175 1.1250 ;
        RECT 5.1975 0.9750 5.5125 1.1250 ;
        RECT 5.0925 0.8250 5.1975 1.1250 ;
        RECT 4.7775 0.9750 5.0925 1.1250 ;
        RECT 4.6725 0.8250 4.7775 1.1250 ;
        RECT 4.3575 0.9750 4.6725 1.1250 ;
        RECT 4.2525 0.8250 4.3575 1.1250 ;
        RECT 3.9375 0.9750 4.2525 1.1250 ;
        RECT 3.8325 0.8250 3.9375 1.1250 ;
        RECT 3.5175 0.9750 3.8325 1.1250 ;
        RECT 3.4125 0.8250 3.5175 1.1250 ;
        RECT 3.0975 0.9750 3.4125 1.1250 ;
        RECT 2.9925 0.8250 3.0975 1.1250 ;
        RECT 2.6775 0.9750 2.9925 1.1250 ;
        RECT 2.5725 0.8250 2.6775 1.1250 ;
        RECT 2.2575 0.9750 2.5725 1.1250 ;
        RECT 2.1525 0.8250 2.2575 1.1250 ;
        RECT 1.8375 0.9750 2.1525 1.1250 ;
        RECT 1.7325 0.8325 1.8375 1.1250 ;
        RECT 1.4175 0.9750 1.7325 1.1250 ;
        RECT 1.3125 0.8250 1.4175 1.1250 ;
        RECT 0.9975 0.9750 1.3125 1.1250 ;
        RECT 0.8925 0.8325 0.9975 1.1250 ;
        RECT 0.5775 0.9750 0.8925 1.1250 ;
        RECT 0.4725 0.8250 0.5775 1.1250 ;
        RECT 0.1575 0.9750 0.4725 1.1250 ;
        RECT 0.0525 0.7875 0.1575 1.1250 ;
        RECT 0.0000 0.9750 0.0525 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 6.7950 0.2100 6.8550 0.2700 ;
        RECT 6.7950 0.8175 6.8550 0.8775 ;
        RECT 6.6900 0.4650 6.7500 0.5250 ;
        RECT 6.5850 0.1275 6.6450 0.1875 ;
        RECT 6.5850 0.7725 6.6450 0.8325 ;
        RECT 6.4800 0.4650 6.5400 0.5250 ;
        RECT 6.3750 0.2700 6.4350 0.3300 ;
        RECT 6.3750 0.8550 6.4350 0.9150 ;
        RECT 6.2700 0.4650 6.3300 0.5250 ;
        RECT 6.1650 0.1275 6.2250 0.1875 ;
        RECT 6.1650 0.6750 6.2250 0.7350 ;
        RECT 6.0600 0.4650 6.1200 0.5250 ;
        RECT 5.9550 0.2700 6.0150 0.3300 ;
        RECT 5.9550 0.8550 6.0150 0.9150 ;
        RECT 5.8500 0.4650 5.9100 0.5250 ;
        RECT 5.7450 0.1275 5.8050 0.1875 ;
        RECT 5.7450 0.6825 5.8050 0.7425 ;
        RECT 5.6400 0.4650 5.7000 0.5250 ;
        RECT 5.5350 0.2700 5.5950 0.3300 ;
        RECT 5.5350 0.8550 5.5950 0.9150 ;
        RECT 5.4300 0.4650 5.4900 0.5250 ;
        RECT 5.3250 0.1275 5.3850 0.1875 ;
        RECT 5.3250 0.6750 5.3850 0.7350 ;
        RECT 5.2200 0.4650 5.2800 0.5250 ;
        RECT 5.1150 0.2700 5.1750 0.3300 ;
        RECT 5.1150 0.8550 5.1750 0.9150 ;
        RECT 5.0100 0.4650 5.0700 0.5250 ;
        RECT 4.9050 0.1275 4.9650 0.1875 ;
        RECT 4.9050 0.6750 4.9650 0.7350 ;
        RECT 4.8000 0.4650 4.8600 0.5250 ;
        RECT 4.6950 0.2700 4.7550 0.3300 ;
        RECT 4.6950 0.8550 4.7550 0.9150 ;
        RECT 4.5900 0.4650 4.6500 0.5250 ;
        RECT 4.4850 0.1275 4.5450 0.1875 ;
        RECT 4.4850 0.6750 4.5450 0.7350 ;
        RECT 4.3800 0.4650 4.4400 0.5250 ;
        RECT 4.2750 0.2700 4.3350 0.3300 ;
        RECT 4.2750 0.8550 4.3350 0.9150 ;
        RECT 4.1700 0.4650 4.2300 0.5250 ;
        RECT 4.0650 0.1275 4.1250 0.1875 ;
        RECT 4.0650 0.6750 4.1250 0.7350 ;
        RECT 3.9600 0.4650 4.0200 0.5250 ;
        RECT 3.8550 0.2700 3.9150 0.3300 ;
        RECT 3.8550 0.8550 3.9150 0.9150 ;
        RECT 3.7500 0.4650 3.8100 0.5250 ;
        RECT 3.6450 0.1275 3.7050 0.1875 ;
        RECT 3.6450 0.6750 3.7050 0.7350 ;
        RECT 3.5400 0.4650 3.6000 0.5250 ;
        RECT 3.4350 0.1575 3.4950 0.2175 ;
        RECT 3.4350 0.8550 3.4950 0.9150 ;
        RECT 3.3300 0.4800 3.3900 0.5400 ;
        RECT 3.2250 0.3000 3.2850 0.3600 ;
        RECT 3.2250 0.6750 3.2850 0.7350 ;
        RECT 3.1200 0.4800 3.1800 0.5400 ;
        RECT 3.0150 0.1575 3.0750 0.2175 ;
        RECT 3.0150 0.8550 3.0750 0.9150 ;
        RECT 2.9100 0.4800 2.9700 0.5400 ;
        RECT 2.8050 0.3000 2.8650 0.3600 ;
        RECT 2.8050 0.6750 2.8650 0.7350 ;
        RECT 2.7000 0.4800 2.7600 0.5400 ;
        RECT 2.5950 0.1575 2.6550 0.2175 ;
        RECT 2.5950 0.8550 2.6550 0.9150 ;
        RECT 2.4900 0.4800 2.5500 0.5400 ;
        RECT 2.3850 0.3000 2.4450 0.3600 ;
        RECT 2.3850 0.6750 2.4450 0.7350 ;
        RECT 2.2800 0.4800 2.3400 0.5400 ;
        RECT 2.1750 0.1575 2.2350 0.2175 ;
        RECT 2.1750 0.8550 2.2350 0.9150 ;
        RECT 2.0700 0.4800 2.1300 0.5400 ;
        RECT 1.9650 0.3000 2.0250 0.3600 ;
        RECT 1.9650 0.6825 2.0250 0.7425 ;
        RECT 1.8600 0.4800 1.9200 0.5400 ;
        RECT 1.7550 0.1575 1.8150 0.2175 ;
        RECT 1.7550 0.8550 1.8150 0.9150 ;
        RECT 1.6500 0.4800 1.7100 0.5400 ;
        RECT 1.5450 0.3000 1.6050 0.3600 ;
        RECT 1.5450 0.6750 1.6050 0.7350 ;
        RECT 1.4400 0.4800 1.5000 0.5400 ;
        RECT 1.3350 0.1575 1.3950 0.2175 ;
        RECT 1.3350 0.8550 1.3950 0.9150 ;
        RECT 1.2300 0.4800 1.2900 0.5400 ;
        RECT 1.1250 0.3000 1.1850 0.3600 ;
        RECT 1.1250 0.6750 1.1850 0.7350 ;
        RECT 1.0200 0.4800 1.0800 0.5400 ;
        RECT 0.9150 0.1575 0.9750 0.2175 ;
        RECT 0.9150 0.8550 0.9750 0.9150 ;
        RECT 0.8100 0.4800 0.8700 0.5400 ;
        RECT 0.1800 0.4800 0.2400 0.5400 ;
        RECT 0.0750 0.1800 0.1350 0.2400 ;
        RECT 0.0750 0.8175 0.1350 0.8775 ;
        RECT 0.7050 0.3000 0.7650 0.3600 ;
        RECT 0.7050 0.6750 0.7650 0.7350 ;
        RECT 0.6000 0.4800 0.6600 0.5400 ;
        RECT 0.4950 0.1575 0.5550 0.2175 ;
        RECT 0.4950 0.8550 0.5550 0.9150 ;
        RECT 0.3900 0.4800 0.4500 0.5400 ;
        RECT 0.2850 0.3000 0.3450 0.3600 ;
        RECT 0.2850 0.7800 0.3450 0.8400 ;
        LAYER M1 ;
        RECT 6.7875 0.1800 6.8625 0.3375 ;
        RECT 3.5325 0.2625 6.7875 0.3375 ;
        RECT 6.5775 0.6675 6.6525 0.8700 ;
        RECT 0.3525 0.6675 6.5775 0.7425 ;
        RECT 3.4575 0.1500 3.5325 0.3375 ;
        RECT 0.1575 0.1500 3.4575 0.2250 ;
        RECT 0.2550 0.3000 3.3825 0.4050 ;
        RECT 0.2775 0.6675 0.3525 0.8700 ;
        RECT 0.0525 0.1500 0.1575 0.2700 ;
        LAYER M2 ;
        RECT 2.8125 0.2925 2.9400 0.4125 ;
        RECT 2.8125 0.6450 2.9400 0.7650 ;
        RECT 2.3100 0.2925 2.4375 0.4125 ;
        RECT 2.3100 0.6450 2.4375 0.7650 ;
    END
END ND2_1100


MACRO ND3_0001
    CLASS CORE ;
    FOREIGN ND3_0001 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.1000 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 1.7475 0.6675 1.8225 0.8700 ;
        RECT 0.1425 0.6675 1.7475 0.7425 ;
        RECT 0.1425 0.3000 0.6000 0.3900 ;
        RECT 0.1125 0.2175 0.1425 0.3900 ;
        RECT 0.1125 0.6675 0.1425 0.8700 ;
        RECT 0.0375 0.2175 0.1125 0.8700 ;
        END
    END ZN
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.9575 0.3675 2.0325 0.6825 ;
        RECT 1.4325 0.4500 1.9575 0.5700 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.9975 0.5625 1.4625 0.6375 ;
        RECT 0.8925 0.4350 0.9975 0.6375 ;
        VIA 0.9450 0.5175 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.5775 0.2625 1.0425 0.3375 ;
        RECT 0.4725 0.2625 0.5775 0.6000 ;
        VIA 0.5250 0.5175 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 2.0325 -0.0750 2.1000 0.0750 ;
        RECT 1.9575 -0.0750 2.0325 0.2475 ;
        RECT 1.6350 -0.0750 1.9575 0.0750 ;
        RECT 1.5150 -0.0750 1.6350 0.2100 ;
        RECT 0.0000 -0.0750 1.5150 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 2.0325 0.9750 2.1000 1.1250 ;
        RECT 1.9575 0.8025 2.0325 1.1250 ;
        RECT 1.6275 0.9750 1.9575 1.1250 ;
        RECT 1.5225 0.8250 1.6275 1.1250 ;
        RECT 1.2075 0.9750 1.5225 1.1250 ;
        RECT 1.1025 0.8250 1.2075 1.1250 ;
        RECT 0.7875 0.9750 1.1025 1.1250 ;
        RECT 0.6825 0.8250 0.7875 1.1250 ;
        RECT 0.3675 0.9750 0.6825 1.1250 ;
        RECT 0.2625 0.8250 0.3675 1.1250 ;
        RECT 0.0000 0.9750 0.2625 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.9650 0.1575 2.0250 0.2175 ;
        RECT 1.9650 0.8325 2.0250 0.8925 ;
        RECT 1.8600 0.4800 1.9200 0.5400 ;
        RECT 1.7550 0.3000 1.8150 0.3600 ;
        RECT 1.7550 0.7725 1.8150 0.8325 ;
        RECT 1.6500 0.4800 1.7100 0.5400 ;
        RECT 1.5450 0.1350 1.6050 0.1950 ;
        RECT 1.5450 0.8550 1.6050 0.9150 ;
        RECT 1.4400 0.4800 1.5000 0.5400 ;
        RECT 1.3350 0.3000 1.3950 0.3600 ;
        RECT 1.3350 0.6750 1.3950 0.7350 ;
        RECT 1.2300 0.4800 1.2900 0.5400 ;
        RECT 1.1250 0.1575 1.1850 0.2175 ;
        RECT 1.1250 0.8550 1.1850 0.9150 ;
        RECT 1.0200 0.4800 1.0800 0.5400 ;
        RECT 0.9150 0.3000 0.9750 0.3600 ;
        RECT 0.9150 0.6750 0.9750 0.7350 ;
        RECT 0.8100 0.4800 0.8700 0.5400 ;
        RECT 0.7050 0.1575 0.7650 0.2175 ;
        RECT 0.7050 0.8550 0.7650 0.9150 ;
        RECT 0.6000 0.4950 0.6600 0.5550 ;
        RECT 0.4950 0.3000 0.5550 0.3600 ;
        RECT 0.4950 0.6750 0.5550 0.7350 ;
        RECT 0.3900 0.4950 0.4500 0.5550 ;
        RECT 0.2850 0.1575 0.3450 0.2175 ;
        RECT 0.2850 0.8550 0.3450 0.9150 ;
        RECT 0.1875 0.4950 0.2475 0.5550 ;
        RECT 0.0750 0.3000 0.1350 0.3600 ;
        RECT 0.0750 0.7800 0.1350 0.8400 ;
        LAYER M1 ;
        RECT 0.8850 0.3000 1.8525 0.3750 ;
        RECT 0.8025 0.4500 1.3125 0.5700 ;
        RECT 0.2550 0.1500 1.2825 0.2250 ;
        RECT 0.1875 0.4650 0.6900 0.5850 ;
    END
END ND3_0001


MACRO ND3_0010
    CLASS CORE ;
    FOREIGN ND3_0010 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.7200 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 1.3125 0.2925 1.4700 0.4125 ;
        RECT 1.3125 0.6300 1.4700 0.7500 ;
        RECT 0.9975 0.2925 1.3125 0.7500 ;
        RECT 0.8400 0.2925 0.9975 0.4125 ;
        RECT 0.8400 0.6300 0.9975 0.7500 ;
        VIA 1.3125 0.3525 VIA12_slot ;
        VIA 1.3125 0.6900 VIA12_slot ;
        VIA 0.9975 0.3525 VIA12_slot ;
        VIA 0.9975 0.6900 VIA12_slot ;
        END
    END ZN
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 6.5325 0.4125 6.6375 0.6825 ;
        RECT 6.4725 0.4125 6.5325 0.5475 ;
        RECT 4.1400 0.4725 6.4725 0.5475 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 2.2575 0.4125 2.3625 0.6000 ;
        RECT 1.8975 0.4125 2.2575 0.4875 ;
        VIA 2.3100 0.5025 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1425 0.4800 1.7400 0.5550 ;
        RECT 0.0675 0.3675 0.1425 0.6825 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 6.4650 -0.0750 6.7200 0.0750 ;
        RECT 6.3450 -0.0750 6.4650 0.1875 ;
        RECT 6.0450 -0.0750 6.3450 0.0750 ;
        RECT 5.9250 -0.0750 6.0450 0.2100 ;
        RECT 5.6250 -0.0750 5.9250 0.0750 ;
        RECT 5.5050 -0.0750 5.6250 0.2100 ;
        RECT 5.2050 -0.0750 5.5050 0.0750 ;
        RECT 5.0850 -0.0750 5.2050 0.2100 ;
        RECT 4.7850 -0.0750 5.0850 0.0750 ;
        RECT 4.6650 -0.0750 4.7850 0.2100 ;
        RECT 4.3650 -0.0750 4.6650 0.0750 ;
        RECT 4.2450 -0.0750 4.3650 0.2100 ;
        RECT 0.0000 -0.0750 4.2450 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 6.6525 0.9750 6.7200 1.1250 ;
        RECT 6.5775 0.7875 6.6525 1.1250 ;
        RECT 6.2475 0.9750 6.5775 1.1250 ;
        RECT 6.1425 0.8250 6.2475 1.1250 ;
        RECT 5.8275 0.9750 6.1425 1.1250 ;
        RECT 5.7225 0.8250 5.8275 1.1250 ;
        RECT 5.4075 0.9750 5.7225 1.1250 ;
        RECT 5.3025 0.8250 5.4075 1.1250 ;
        RECT 4.9875 0.9750 5.3025 1.1250 ;
        RECT 4.8825 0.8250 4.9875 1.1250 ;
        RECT 4.5675 0.9750 4.8825 1.1250 ;
        RECT 4.4625 0.8250 4.5675 1.1250 ;
        RECT 4.1550 0.9750 4.4625 1.1250 ;
        RECT 4.0350 0.8250 4.1550 1.1250 ;
        RECT 3.9450 0.9750 4.0350 1.1250 ;
        RECT 3.8250 0.8250 3.9450 1.1250 ;
        RECT 3.5250 0.9750 3.8250 1.1250 ;
        RECT 3.4050 0.8250 3.5250 1.1250 ;
        RECT 3.0975 0.9750 3.4050 1.1250 ;
        RECT 2.9925 0.8250 3.0975 1.1250 ;
        RECT 2.6775 0.9750 2.9925 1.1250 ;
        RECT 2.5725 0.8250 2.6775 1.1250 ;
        RECT 2.2575 0.9750 2.5725 1.1250 ;
        RECT 2.1525 0.8250 2.2575 1.1250 ;
        RECT 1.8375 0.9750 2.1525 1.1250 ;
        RECT 1.7325 0.8250 1.8375 1.1250 ;
        RECT 1.4175 0.9750 1.7325 1.1250 ;
        RECT 1.3125 0.8250 1.4175 1.1250 ;
        RECT 0.9975 0.9750 1.3125 1.1250 ;
        RECT 0.8925 0.8250 0.9975 1.1250 ;
        RECT 0.5775 0.9750 0.8925 1.1250 ;
        RECT 0.4725 0.8250 0.5775 1.1250 ;
        RECT 0.1425 0.9750 0.4725 1.1250 ;
        RECT 0.0675 0.8025 0.1425 1.1250 ;
        RECT 0.0000 0.9750 0.0675 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 6.5850 0.2100 6.6450 0.2700 ;
        RECT 6.5850 0.8325 6.6450 0.8925 ;
        RECT 6.4800 0.4800 6.5400 0.5400 ;
        RECT 6.3750 0.1275 6.4350 0.1875 ;
        RECT 6.3750 0.8175 6.4350 0.8775 ;
        RECT 6.2700 0.4800 6.3300 0.5400 ;
        RECT 6.1650 0.3000 6.2250 0.3600 ;
        RECT 6.1650 0.8550 6.2250 0.9150 ;
        RECT 6.0600 0.4800 6.1200 0.5400 ;
        RECT 5.9550 0.1350 6.0150 0.1950 ;
        RECT 5.9550 0.8175 6.0150 0.8775 ;
        RECT 5.8500 0.4800 5.9100 0.5400 ;
        RECT 5.7450 0.3000 5.8050 0.3600 ;
        RECT 5.7450 0.8550 5.8050 0.9150 ;
        RECT 5.6400 0.4800 5.7000 0.5400 ;
        RECT 5.5350 0.1350 5.5950 0.1950 ;
        RECT 5.5350 0.8175 5.5950 0.8775 ;
        RECT 5.4300 0.4800 5.4900 0.5400 ;
        RECT 5.3250 0.3000 5.3850 0.3600 ;
        RECT 5.3250 0.8550 5.3850 0.9150 ;
        RECT 5.2200 0.4800 5.2800 0.5400 ;
        RECT 5.1150 0.1350 5.1750 0.1950 ;
        RECT 5.1150 0.8175 5.1750 0.8775 ;
        RECT 5.0100 0.4800 5.0700 0.5400 ;
        RECT 4.9050 0.3000 4.9650 0.3600 ;
        RECT 4.9050 0.8550 4.9650 0.9150 ;
        RECT 4.8000 0.4800 4.8600 0.5400 ;
        RECT 4.6950 0.1350 4.7550 0.1950 ;
        RECT 4.6950 0.6600 4.7550 0.7200 ;
        RECT 4.5900 0.4800 4.6500 0.5400 ;
        RECT 4.4850 0.3000 4.5450 0.3600 ;
        RECT 4.4850 0.8550 4.5450 0.9150 ;
        RECT 4.3800 0.4800 4.4400 0.5400 ;
        RECT 4.2750 0.1350 4.3350 0.1950 ;
        RECT 4.2750 0.6600 4.3350 0.7200 ;
        RECT 4.1700 0.4800 4.2300 0.5400 ;
        RECT 4.0650 0.3000 4.1250 0.3600 ;
        RECT 4.0650 0.8325 4.1250 0.8925 ;
        RECT 3.8550 0.1575 3.9150 0.2175 ;
        RECT 3.8550 0.8325 3.9150 0.8925 ;
        RECT 3.7500 0.4800 3.8100 0.5400 ;
        RECT 3.6450 0.3000 3.7050 0.3600 ;
        RECT 3.6450 0.8175 3.7050 0.8775 ;
        RECT 3.5400 0.4800 3.6000 0.5400 ;
        RECT 3.4350 0.1575 3.4950 0.2175 ;
        RECT 3.4350 0.8325 3.4950 0.8925 ;
        RECT 3.3300 0.4800 3.3900 0.5400 ;
        RECT 3.2250 0.3000 3.2850 0.3600 ;
        RECT 3.2250 0.8175 3.2850 0.8775 ;
        RECT 3.1200 0.4800 3.1800 0.5400 ;
        RECT 3.0150 0.1575 3.0750 0.2175 ;
        RECT 3.0150 0.8550 3.0750 0.9150 ;
        RECT 2.9100 0.4800 2.9700 0.5400 ;
        RECT 2.8050 0.3000 2.8650 0.3600 ;
        RECT 2.8050 0.6600 2.8650 0.7200 ;
        RECT 2.7000 0.4800 2.7600 0.5400 ;
        RECT 2.5950 0.1575 2.6550 0.2175 ;
        RECT 2.5950 0.8550 2.6550 0.9150 ;
        RECT 2.4900 0.4800 2.5500 0.5400 ;
        RECT 2.3850 0.3000 2.4450 0.3600 ;
        RECT 2.3850 0.6600 2.4450 0.7200 ;
        RECT 2.2800 0.4800 2.3400 0.5400 ;
        RECT 2.1750 0.1575 2.2350 0.2175 ;
        RECT 2.1750 0.8550 2.2350 0.9150 ;
        RECT 2.0700 0.4800 2.1300 0.5400 ;
        RECT 1.9650 0.3000 2.0250 0.3600 ;
        RECT 1.9650 0.6600 2.0250 0.7200 ;
        RECT 1.8675 0.4800 1.9275 0.5400 ;
        RECT 1.7550 0.1575 1.8150 0.2175 ;
        RECT 1.7550 0.8550 1.8150 0.9150 ;
        RECT 1.6500 0.4800 1.7100 0.5400 ;
        RECT 1.5450 0.3000 1.6050 0.3600 ;
        RECT 1.5450 0.6600 1.6050 0.7200 ;
        RECT 1.4400 0.4800 1.5000 0.5400 ;
        RECT 1.3350 0.1575 1.3950 0.2175 ;
        RECT 1.3350 0.8550 1.3950 0.9150 ;
        RECT 1.2300 0.4800 1.2900 0.5400 ;
        RECT 1.1250 0.3000 1.1850 0.3600 ;
        RECT 1.1250 0.6600 1.1850 0.7200 ;
        RECT 1.0200 0.4800 1.0800 0.5400 ;
        RECT 0.9150 0.1575 0.9750 0.2175 ;
        RECT 0.9150 0.8550 0.9750 0.9150 ;
        RECT 0.8100 0.4800 0.8700 0.5400 ;
        RECT 0.7050 0.3000 0.7650 0.3600 ;
        RECT 0.7050 0.6600 0.7650 0.7200 ;
        RECT 0.6000 0.4800 0.6600 0.5400 ;
        RECT 0.4950 0.1575 0.5550 0.2175 ;
        RECT 0.4950 0.8550 0.5550 0.9150 ;
        RECT 0.3900 0.4800 0.4500 0.5400 ;
        RECT 0.2850 0.3000 0.3450 0.3600 ;
        RECT 0.2850 0.6600 0.3450 0.7200 ;
        RECT 0.1800 0.4800 0.2400 0.5400 ;
        RECT 0.0750 0.1725 0.1350 0.2325 ;
        RECT 0.0750 0.8325 0.1350 0.8925 ;
        LAYER M1 ;
        RECT 6.5775 0.1800 6.6525 0.3375 ;
        RECT 6.3975 0.2625 6.5775 0.3375 ;
        RECT 6.3525 0.6300 6.4575 0.9000 ;
        RECT 6.3225 0.2625 6.3975 0.3750 ;
        RECT 6.0375 0.6300 6.3525 0.7500 ;
        RECT 1.9350 0.3000 6.3225 0.3750 ;
        RECT 5.9325 0.6300 6.0375 0.9000 ;
        RECT 5.6175 0.6300 5.9325 0.7500 ;
        RECT 5.5125 0.6300 5.6175 0.9000 ;
        RECT 5.1975 0.6300 5.5125 0.7500 ;
        RECT 5.0925 0.6300 5.1975 0.9000 ;
        RECT 3.7275 0.6300 5.0925 0.7500 ;
        RECT 0.1575 0.1500 3.9600 0.2250 ;
        RECT 1.9650 0.4500 3.8625 0.5550 ;
        RECT 3.6225 0.6300 3.7275 0.9000 ;
        RECT 3.3075 0.6300 3.6225 0.7500 ;
        RECT 3.2025 0.6300 3.3075 0.9000 ;
        RECT 2.0475 0.6300 3.2025 0.7500 ;
        RECT 1.8075 0.6375 2.0475 0.7500 ;
        RECT 1.8450 0.4500 1.9650 0.5625 ;
        RECT 0.2775 0.6300 1.8075 0.7500 ;
        RECT 0.2550 0.3000 1.6500 0.4050 ;
        RECT 0.0525 0.1500 0.1575 0.2550 ;
        LAYER M2 ;
        RECT 1.3425 0.2925 1.4700 0.4125 ;
        RECT 1.3425 0.6300 1.4700 0.7500 ;
        RECT 0.8400 0.2925 0.9675 0.4125 ;
        RECT 0.8400 0.6300 0.9675 0.7500 ;
    END
END ND3_0010


MACRO ND3_0011
    CLASS CORE ;
    FOREIGN ND3_0011 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.4700 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 0.8625 0.1125 0.9375 0.7800 ;
        RECT 0.4425 0.1125 0.8625 0.1875 ;
        RECT 0.7725 0.7050 0.8625 0.7800 ;
        VIA 0.9000 0.2025 VIA12_square ;
        VIA 0.8550 0.7425 VIA12_square ;
        END
    END ZN
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.2225 0.3150 1.3275 0.5700 ;
        RECT 0.2475 0.3150 1.2225 0.3900 ;
        RECT 0.1425 0.3150 0.2475 0.5700 ;
        RECT 0.0675 0.3150 0.1425 0.6825 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.0125 0.4650 1.1175 0.9375 ;
        RECT 0.4575 0.8625 1.0125 0.9375 ;
        RECT 0.3825 0.4650 0.4575 0.9375 ;
        VIA 1.0650 0.5475 VIA12_square ;
        VIA 0.4200 0.5775 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.6825 0.2625 0.7875 0.6300 ;
        RECT 0.2175 0.2625 0.6825 0.3375 ;
        VIA 0.7350 0.5475 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.4175 -0.0750 1.4700 0.0750 ;
        RECT 1.3125 -0.0750 1.4175 0.2400 ;
        RECT 0.1575 -0.0750 1.3125 0.0750 ;
        RECT 0.0525 -0.0750 0.1575 0.2400 ;
        RECT 0.0000 -0.0750 0.0525 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.4175 0.9750 1.4700 1.1250 ;
        RECT 1.3125 0.6450 1.4175 1.1250 ;
        RECT 1.0050 0.9750 1.3125 1.1250 ;
        RECT 0.8850 0.8625 1.0050 1.1250 ;
        RECT 0.5850 0.9750 0.8850 1.1250 ;
        RECT 0.4650 0.8625 0.5850 1.1250 ;
        RECT 0.1425 0.9750 0.4650 1.1250 ;
        RECT 0.0675 0.7875 0.1425 1.1250 ;
        RECT 0.0000 0.9750 0.0675 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.3350 0.1575 1.3950 0.2175 ;
        RECT 1.3350 0.6675 1.3950 0.7275 ;
        RECT 1.3350 0.8325 1.3950 0.8925 ;
        RECT 1.2300 0.4800 1.2900 0.5400 ;
        RECT 1.1250 0.7125 1.1850 0.7725 ;
        RECT 1.0200 0.4800 1.0800 0.5400 ;
        RECT 0.9150 0.8625 0.9750 0.9225 ;
        RECT 0.8100 0.4950 0.8700 0.5550 ;
        RECT 0.7050 0.1650 0.7650 0.2250 ;
        RECT 0.7050 0.7125 0.7650 0.7725 ;
        RECT 0.6000 0.4950 0.6600 0.5550 ;
        RECT 0.4950 0.8625 0.5550 0.9225 ;
        RECT 0.3900 0.4800 0.4500 0.5400 ;
        RECT 0.2850 0.7125 0.3450 0.7725 ;
        RECT 0.1800 0.4800 0.2400 0.5400 ;
        RECT 0.0750 0.1575 0.1350 0.2175 ;
        RECT 0.0750 0.8175 0.1350 0.8775 ;
        LAYER M1 ;
        RECT 1.1025 0.7050 1.2375 0.8100 ;
        RECT 0.6750 0.1500 1.2000 0.2400 ;
        RECT 0.9525 0.4650 1.1475 0.6300 ;
        RECT 0.2550 0.7050 1.1025 0.7800 ;
        RECT 0.5925 0.4650 0.8775 0.6300 ;
        RECT 0.3225 0.4650 0.5175 0.6300 ;
    END
END ND3_0011


MACRO ND3_0100
    CLASS CORE ;
    FOREIGN ND3_0100 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.4600 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 1.1025 0.2925 1.2600 0.4125 ;
        RECT 1.1025 0.6300 1.2600 0.7500 ;
        RECT 0.7875 0.2925 1.1025 0.7500 ;
        RECT 0.6300 0.2925 0.7875 0.4125 ;
        RECT 0.6300 0.6300 0.7875 0.7500 ;
        VIA 1.1025 0.3525 VIA12_slot ;
        VIA 1.1025 0.6900 VIA12_slot ;
        VIA 0.7875 0.3525 VIA12_slot ;
        VIA 0.7875 0.6900 VIA12_slot ;
        END
    END ZN
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 3.8700 0.4275 3.9750 0.6375 ;
        RECT 3.4050 0.5625 3.8700 0.6375 ;
        VIA 3.9225 0.5100 VIA12_square ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 2.3625 0.4125 2.4675 0.6000 ;
        RECT 1.8975 0.4125 2.3625 0.4875 ;
        VIA 2.4150 0.5025 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1425 0.4800 1.7400 0.5550 ;
        RECT 0.0675 0.3675 0.1425 0.6825 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 5.2050 -0.0750 5.4600 0.0750 ;
        RECT 5.0850 -0.0750 5.2050 0.2100 ;
        RECT 4.7850 -0.0750 5.0850 0.0750 ;
        RECT 4.6650 -0.0750 4.7850 0.2100 ;
        RECT 4.3650 -0.0750 4.6650 0.0750 ;
        RECT 4.2450 -0.0750 4.3650 0.2100 ;
        RECT 3.9450 -0.0750 4.2450 0.0750 ;
        RECT 3.8250 -0.0750 3.9450 0.2100 ;
        RECT 0.0000 -0.0750 3.8250 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 5.4075 0.9750 5.4600 1.1250 ;
        RECT 5.3025 0.6450 5.4075 1.1250 ;
        RECT 4.9875 0.9750 5.3025 1.1250 ;
        RECT 4.8825 0.8250 4.9875 1.1250 ;
        RECT 4.5675 0.9750 4.8825 1.1250 ;
        RECT 4.4625 0.8250 4.5675 1.1250 ;
        RECT 4.1475 0.9750 4.4625 1.1250 ;
        RECT 4.0425 0.8250 4.1475 1.1250 ;
        RECT 3.7350 0.9750 4.0425 1.1250 ;
        RECT 3.6150 0.8250 3.7350 1.1250 ;
        RECT 3.5250 0.9750 3.6150 1.1250 ;
        RECT 3.4050 0.8250 3.5250 1.1250 ;
        RECT 3.0975 0.9750 3.4050 1.1250 ;
        RECT 2.9925 0.8250 3.0975 1.1250 ;
        RECT 2.6775 0.9750 2.9925 1.1250 ;
        RECT 2.5725 0.8250 2.6775 1.1250 ;
        RECT 2.2575 0.9750 2.5725 1.1250 ;
        RECT 2.1525 0.8250 2.2575 1.1250 ;
        RECT 1.8375 0.9750 2.1525 1.1250 ;
        RECT 1.7325 0.8250 1.8375 1.1250 ;
        RECT 1.4175 0.9750 1.7325 1.1250 ;
        RECT 1.3125 0.8250 1.4175 1.1250 ;
        RECT 0.9975 0.9750 1.3125 1.1250 ;
        RECT 0.8925 0.8250 0.9975 1.1250 ;
        RECT 0.5775 0.9750 0.8925 1.1250 ;
        RECT 0.4725 0.8250 0.5775 1.1250 ;
        RECT 0.1425 0.9750 0.4725 1.1250 ;
        RECT 0.0675 0.8025 0.1425 1.1250 ;
        RECT 0.0000 0.9750 0.0675 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 5.3250 0.2100 5.3850 0.2700 ;
        RECT 5.3250 0.6675 5.3850 0.7275 ;
        RECT 5.3250 0.8325 5.3850 0.8925 ;
        RECT 5.2200 0.4800 5.2800 0.5400 ;
        RECT 5.1150 0.1350 5.1750 0.1950 ;
        RECT 5.1150 0.6600 5.1750 0.7200 ;
        RECT 5.0100 0.4800 5.0700 0.5400 ;
        RECT 4.9050 0.3000 4.9650 0.3600 ;
        RECT 4.9050 0.8550 4.9650 0.9150 ;
        RECT 4.8000 0.4800 4.8600 0.5400 ;
        RECT 4.6950 0.1350 4.7550 0.1950 ;
        RECT 4.6950 0.6600 4.7550 0.7200 ;
        RECT 4.5900 0.4800 4.6500 0.5400 ;
        RECT 4.4850 0.3000 4.5450 0.3600 ;
        RECT 4.4850 0.8550 4.5450 0.9150 ;
        RECT 4.3800 0.4800 4.4400 0.5400 ;
        RECT 4.2750 0.1350 4.3350 0.1950 ;
        RECT 4.2750 0.6600 4.3350 0.7200 ;
        RECT 4.1700 0.4800 4.2300 0.5400 ;
        RECT 4.0650 0.3000 4.1250 0.3600 ;
        RECT 4.0650 0.8550 4.1250 0.9150 ;
        RECT 3.9600 0.4800 4.0200 0.5400 ;
        RECT 3.8550 0.1350 3.9150 0.1950 ;
        RECT 3.8550 0.6600 3.9150 0.7200 ;
        RECT 3.7500 0.4800 3.8100 0.5400 ;
        RECT 3.6450 0.3000 3.7050 0.3600 ;
        RECT 3.6450 0.8325 3.7050 0.8925 ;
        RECT 3.4350 0.1575 3.4950 0.2175 ;
        RECT 3.4350 0.8325 3.4950 0.8925 ;
        RECT 3.3300 0.4800 3.3900 0.5400 ;
        RECT 3.2250 0.3000 3.2850 0.3600 ;
        RECT 3.2250 0.6600 3.2850 0.7200 ;
        RECT 3.1200 0.4800 3.1800 0.5400 ;
        RECT 3.0150 0.1575 3.0750 0.2175 ;
        RECT 3.0150 0.8550 3.0750 0.9150 ;
        RECT 2.9100 0.4800 2.9700 0.5400 ;
        RECT 2.8050 0.3000 2.8650 0.3600 ;
        RECT 2.8050 0.6600 2.8650 0.7200 ;
        RECT 2.7000 0.4800 2.7600 0.5400 ;
        RECT 2.5950 0.1575 2.6550 0.2175 ;
        RECT 2.5950 0.8550 2.6550 0.9150 ;
        RECT 2.4900 0.4800 2.5500 0.5400 ;
        RECT 2.3850 0.3000 2.4450 0.3600 ;
        RECT 2.3850 0.6600 2.4450 0.7200 ;
        RECT 2.2800 0.4800 2.3400 0.5400 ;
        RECT 2.1750 0.1575 2.2350 0.2175 ;
        RECT 2.1750 0.8550 2.2350 0.9150 ;
        RECT 2.0700 0.4800 2.1300 0.5400 ;
        RECT 1.9650 0.3000 2.0250 0.3600 ;
        RECT 1.9650 0.6600 2.0250 0.7200 ;
        RECT 1.8600 0.4800 1.9200 0.5400 ;
        RECT 1.7550 0.1575 1.8150 0.2175 ;
        RECT 1.7550 0.8550 1.8150 0.9150 ;
        RECT 1.6500 0.4800 1.7100 0.5400 ;
        RECT 1.5450 0.3000 1.6050 0.3600 ;
        RECT 1.5450 0.6600 1.6050 0.7200 ;
        RECT 1.4400 0.4800 1.5000 0.5400 ;
        RECT 1.3350 0.1575 1.3950 0.2175 ;
        RECT 1.3350 0.8550 1.3950 0.9150 ;
        RECT 1.2300 0.4800 1.2900 0.5400 ;
        RECT 1.1250 0.3000 1.1850 0.3600 ;
        RECT 1.1250 0.6600 1.1850 0.7200 ;
        RECT 1.0200 0.4800 1.0800 0.5400 ;
        RECT 0.9150 0.1575 0.9750 0.2175 ;
        RECT 0.9150 0.8550 0.9750 0.9150 ;
        RECT 0.8100 0.4800 0.8700 0.5400 ;
        RECT 0.7050 0.3000 0.7650 0.3600 ;
        RECT 0.7050 0.6600 0.7650 0.7200 ;
        RECT 0.6000 0.4800 0.6600 0.5400 ;
        RECT 0.4950 0.1575 0.5550 0.2175 ;
        RECT 0.4950 0.8550 0.5550 0.9150 ;
        RECT 0.3900 0.4800 0.4500 0.5400 ;
        RECT 0.2850 0.3000 0.3450 0.3600 ;
        RECT 0.2850 0.6600 0.3450 0.7200 ;
        RECT 0.1800 0.4800 0.2400 0.5400 ;
        RECT 0.0750 0.1725 0.1350 0.2325 ;
        RECT 0.0750 0.8325 0.1350 0.8925 ;
        LAYER M1 ;
        RECT 5.3175 0.1800 5.3925 0.3750 ;
        RECT 3.7200 0.4725 5.3250 0.5475 ;
        RECT 1.9350 0.3000 5.3175 0.3750 ;
        RECT 2.0475 0.6300 5.1825 0.7500 ;
        RECT 0.1575 0.1500 3.5400 0.2250 ;
        RECT 1.9650 0.4500 3.4425 0.5550 ;
        RECT 1.8075 0.6450 2.0475 0.7500 ;
        RECT 1.8600 0.4500 1.9650 0.5700 ;
        RECT 0.2775 0.6300 1.8075 0.7500 ;
        RECT 0.2550 0.3000 1.6500 0.4050 ;
        RECT 0.0525 0.1500 0.1575 0.2550 ;
        LAYER M2 ;
        RECT 1.1325 0.2925 1.2600 0.4125 ;
        RECT 1.1325 0.6300 1.2600 0.7500 ;
        RECT 0.6300 0.2925 0.7575 0.4125 ;
        RECT 0.6300 0.6300 0.7575 0.7500 ;
    END
END ND3_0100


MACRO ND3_0111
    CLASS CORE ;
    FOREIGN ND3_0111 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.9400 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 0.3675 0.2700 0.6825 0.7875 ;
        VIA 0.5250 0.3525 VIA12_slot ;
        VIA 0.5250 0.7050 VIA12_slot ;
        END
    END ZN
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 2.2275 0.4125 2.5275 0.4875 ;
        RECT 2.1525 0.4125 2.2275 0.5775 ;
        RECT 1.9875 0.4125 2.1525 0.4875 ;
        VIA 2.1900 0.4950 VIA12_square ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.5375 0.4125 1.6125 0.5775 ;
        RECT 1.0725 0.4125 1.5375 0.4875 ;
        VIA 1.5750 0.4950 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1425 0.4800 0.9000 0.5850 ;
        RECT 0.0675 0.3675 0.1425 0.6825 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 2.6850 -0.0750 2.9400 0.0750 ;
        RECT 2.5650 -0.0750 2.6850 0.2100 ;
        RECT 2.2650 -0.0750 2.5650 0.0750 ;
        RECT 2.1450 -0.0750 2.2650 0.2100 ;
        RECT 0.0000 -0.0750 2.1450 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 2.8725 0.9750 2.9400 1.1250 ;
        RECT 2.7975 0.8025 2.8725 1.1250 ;
        RECT 2.4675 0.9750 2.7975 1.1250 ;
        RECT 2.3625 0.8250 2.4675 1.1250 ;
        RECT 2.0550 0.9750 2.3625 1.1250 ;
        RECT 1.9350 0.8175 2.0550 1.1250 ;
        RECT 1.8450 0.9750 1.9350 1.1250 ;
        RECT 1.7250 0.8175 1.8450 1.1250 ;
        RECT 1.4175 0.9750 1.7250 1.1250 ;
        RECT 1.3125 0.8250 1.4175 1.1250 ;
        RECT 0.9975 0.9750 1.3125 1.1250 ;
        RECT 0.8925 0.8250 0.9975 1.1250 ;
        RECT 0.5775 0.9750 0.8925 1.1250 ;
        RECT 0.4725 0.8250 0.5775 1.1250 ;
        RECT 0.1650 0.9750 0.4725 1.1250 ;
        RECT 0.0450 0.8250 0.1650 1.1250 ;
        RECT 0.0000 0.9750 0.0450 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 2.8050 0.2100 2.8650 0.2700 ;
        RECT 2.8050 0.8325 2.8650 0.8925 ;
        RECT 2.7000 0.4800 2.7600 0.5400 ;
        RECT 2.5950 0.1350 2.6550 0.1950 ;
        RECT 2.5950 0.7725 2.6550 0.8325 ;
        RECT 2.4900 0.4800 2.5500 0.5400 ;
        RECT 2.3850 0.3000 2.4450 0.3600 ;
        RECT 2.3850 0.8550 2.4450 0.9150 ;
        RECT 2.2800 0.4800 2.3400 0.5400 ;
        RECT 2.1750 0.1350 2.2350 0.1950 ;
        RECT 2.1750 0.6750 2.2350 0.7350 ;
        RECT 2.0700 0.4800 2.1300 0.5400 ;
        RECT 1.9650 0.3000 2.0250 0.3600 ;
        RECT 1.9650 0.8325 2.0250 0.8925 ;
        RECT 1.7550 0.1575 1.8150 0.2175 ;
        RECT 1.7550 0.8325 1.8150 0.8925 ;
        RECT 1.6500 0.4800 1.7100 0.5400 ;
        RECT 1.5450 0.3000 1.6050 0.3600 ;
        RECT 1.5450 0.6750 1.6050 0.7350 ;
        RECT 1.4400 0.4800 1.5000 0.5400 ;
        RECT 1.3350 0.1575 1.3950 0.2175 ;
        RECT 1.3350 0.8550 1.3950 0.9150 ;
        RECT 1.2300 0.4800 1.2900 0.5400 ;
        RECT 1.1250 0.3000 1.1850 0.3600 ;
        RECT 1.1250 0.6750 1.1850 0.7350 ;
        RECT 1.0200 0.4800 1.0800 0.5400 ;
        RECT 0.9150 0.1575 0.9750 0.2175 ;
        RECT 0.9150 0.8550 0.9750 0.9150 ;
        RECT 0.8100 0.4800 0.8700 0.5400 ;
        RECT 0.7050 0.3000 0.7650 0.3600 ;
        RECT 0.7050 0.6750 0.7650 0.7350 ;
        RECT 0.6000 0.4800 0.6600 0.5400 ;
        RECT 0.4950 0.1575 0.5550 0.2175 ;
        RECT 0.4950 0.8550 0.5550 0.9150 ;
        RECT 0.3900 0.4800 0.4500 0.5400 ;
        RECT 0.2850 0.3000 0.3450 0.3600 ;
        RECT 0.2850 0.7800 0.3450 0.8400 ;
        RECT 0.1800 0.4800 0.2400 0.5400 ;
        RECT 0.0750 0.1575 0.1350 0.2175 ;
        RECT 0.0750 0.8325 0.1350 0.8925 ;
        LAYER M1 ;
        RECT 2.7975 0.1800 2.8725 0.3750 ;
        RECT 1.0950 0.3000 2.7975 0.3750 ;
        RECT 2.0625 0.4500 2.7675 0.5700 ;
        RECT 2.5875 0.6675 2.6625 0.8700 ;
        RECT 0.3525 0.6675 2.5875 0.7425 ;
        RECT 0.1575 0.1500 1.8600 0.2250 ;
        RECT 1.0125 0.4500 1.7175 0.5700 ;
        RECT 0.2550 0.3000 0.8100 0.4050 ;
        RECT 0.2775 0.6675 0.3525 0.8700 ;
        RECT 0.0450 0.1500 0.1575 0.2550 ;
    END
END ND3_0111


MACRO ND3_1000
    CLASS CORE ;
    FOREIGN ND3_1000 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.8400 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.7275 0.1500 0.8025 0.9000 ;
        RECT 0.6975 0.1500 0.7275 0.2700 ;
        RECT 0.6825 0.6675 0.7275 0.9000 ;
        RECT 0.3675 0.6675 0.6825 0.7425 ;
        RECT 0.2625 0.6675 0.3675 0.9000 ;
        END
    END ZN
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1425 0.4350 0.2475 0.5550 ;
        RECT 0.0675 0.3675 0.1425 0.6825 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.4725 0.8625 0.7725 0.9375 ;
        RECT 0.3675 0.4275 0.4725 0.9375 ;
        RECT 0.2025 0.8625 0.3675 0.9375 ;
        VIA 0.4200 0.5100 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.3075 0.2625 0.7725 0.3375 ;
        VIA 0.5850 0.3000 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.1650 -0.0750 0.8400 0.0750 ;
        RECT 0.0450 -0.0750 0.1650 0.2475 ;
        RECT 0.0000 -0.0750 0.0450 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.5775 0.9750 0.8400 1.1250 ;
        RECT 0.4725 0.8475 0.5775 1.1250 ;
        RECT 0.1650 0.9750 0.4725 1.1250 ;
        RECT 0.0450 0.8025 0.1650 1.1250 ;
        RECT 0.0000 0.9750 0.0450 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 0.7050 0.1800 0.7650 0.2400 ;
        RECT 0.7050 0.8175 0.7650 0.8775 ;
        RECT 0.5925 0.4650 0.6525 0.5250 ;
        RECT 0.4950 0.8700 0.5550 0.9300 ;
        RECT 0.3900 0.4650 0.4500 0.5250 ;
        RECT 0.2850 0.8175 0.3450 0.8775 ;
        RECT 0.1800 0.4650 0.2400 0.5250 ;
        RECT 0.0750 0.1575 0.1350 0.2175 ;
        RECT 0.0750 0.8325 0.1350 0.8925 ;
        LAYER M1 ;
        RECT 0.6225 0.4350 0.6525 0.5925 ;
        RECT 0.5400 0.2175 0.6225 0.5925 ;
        RECT 0.3225 0.3375 0.4650 0.5925 ;
    END
END ND3_1000


MACRO ND3_1010
    CLASS CORE ;
    FOREIGN ND3_1010 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.8400 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.7275 0.1575 0.8025 0.8325 ;
        RECT 0.6975 0.1575 0.7275 0.2775 ;
        RECT 0.6975 0.6675 0.7275 0.8325 ;
        RECT 0.2550 0.6675 0.6975 0.7425 ;
        END
    END ZN
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1425 0.4350 0.2475 0.5550 ;
        RECT 0.0675 0.3675 0.1425 0.6825 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.3450 0.2175 0.4500 0.5925 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.6225 0.4350 0.6525 0.5925 ;
        RECT 0.5400 0.2175 0.6225 0.5925 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.1650 -0.0750 0.8400 0.0750 ;
        RECT 0.0450 -0.0750 0.1650 0.2475 ;
        RECT 0.0000 -0.0750 0.0450 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.5775 0.9750 0.8400 1.1250 ;
        RECT 0.4725 0.8475 0.5775 1.1250 ;
        RECT 0.1650 0.9750 0.4725 1.1250 ;
        RECT 0.0450 0.8025 0.1650 1.1250 ;
        RECT 0.0000 0.9750 0.0450 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 0.7050 0.1875 0.7650 0.2475 ;
        RECT 0.7050 0.7200 0.7650 0.7800 ;
        RECT 0.5925 0.4650 0.6525 0.5250 ;
        RECT 0.4950 0.8700 0.5550 0.9300 ;
        RECT 0.3900 0.4650 0.4500 0.5250 ;
        RECT 0.2850 0.6750 0.3450 0.7350 ;
        RECT 0.1800 0.4650 0.2400 0.5250 ;
        RECT 0.0750 0.1575 0.1350 0.2175 ;
        RECT 0.0750 0.8325 0.1350 0.8925 ;
    END
END ND3_1010


MACRO ND4_0001
    CLASS CORE ;
    FOREIGN ND4_0001 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.7300 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 2.5725 0.6675 2.6775 0.7875 ;
        RECT 0.1425 0.6675 2.5725 0.7425 ;
        RECT 0.1425 0.3000 0.6000 0.3900 ;
        RECT 0.1125 0.2175 0.1425 0.3900 ;
        RECT 0.1125 0.6675 0.1425 0.8700 ;
        RECT 0.0375 0.2175 0.1125 0.8700 ;
        END
    END ZN
    PIN A4
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 2.1750 0.2625 2.2800 0.6000 ;
        RECT 1.7100 0.2625 2.1750 0.3375 ;
        VIA 2.2275 0.5100 VIA12_square ;
        END
    END A4
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.7325 0.4125 1.8375 0.6300 ;
        RECT 1.2675 0.4125 1.7325 0.4875 ;
        VIA 1.7850 0.5325 VIA12_square ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.9975 0.5625 1.4625 0.6375 ;
        RECT 0.8925 0.4350 0.9975 0.6375 ;
        VIA 0.9450 0.5175 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.5775 0.2625 1.0425 0.3375 ;
        RECT 0.4725 0.2625 0.5775 0.6000 ;
        VIA 0.5250 0.5175 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 2.6625 -0.0750 2.7300 0.0750 ;
        RECT 2.5875 -0.0750 2.6625 0.2550 ;
        RECT 2.2575 -0.0750 2.5875 0.0750 ;
        RECT 2.1525 -0.0750 2.2575 0.2250 ;
        RECT 0.0000 -0.0750 2.1525 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 2.4675 0.9750 2.7300 1.1250 ;
        RECT 2.3625 0.8325 2.4675 1.1250 ;
        RECT 2.0475 0.9750 2.3625 1.1250 ;
        RECT 1.9425 0.8325 2.0475 1.1250 ;
        RECT 1.6350 0.9750 1.9425 1.1250 ;
        RECT 1.5150 0.8325 1.6350 1.1250 ;
        RECT 1.2075 0.9750 1.5150 1.1250 ;
        RECT 1.1025 0.8250 1.2075 1.1250 ;
        RECT 0.7875 0.9750 1.1025 1.1250 ;
        RECT 0.6825 0.8250 0.7875 1.1250 ;
        RECT 0.3675 0.9750 0.6825 1.1250 ;
        RECT 0.2625 0.8250 0.3675 1.1250 ;
        RECT 0.0000 0.9750 0.2625 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 2.5950 0.1575 2.6550 0.2175 ;
        RECT 2.5950 0.6975 2.6550 0.7575 ;
        RECT 2.4900 0.4800 2.5500 0.5400 ;
        RECT 2.3850 0.2175 2.4450 0.2775 ;
        RECT 2.3850 0.8550 2.4450 0.9150 ;
        RECT 2.2800 0.4800 2.3400 0.5400 ;
        RECT 2.1750 0.1425 2.2350 0.2025 ;
        RECT 2.1750 0.6750 2.2350 0.7350 ;
        RECT 2.0700 0.4800 2.1300 0.5400 ;
        RECT 1.9650 0.2400 2.0250 0.3000 ;
        RECT 1.9650 0.8550 2.0250 0.9150 ;
        RECT 1.8600 0.4875 1.9200 0.5475 ;
        RECT 1.7550 0.3075 1.8150 0.3675 ;
        RECT 1.7550 0.6750 1.8150 0.7350 ;
        RECT 1.6500 0.4800 1.7100 0.5400 ;
        RECT 1.5450 0.1575 1.6050 0.2175 ;
        RECT 1.5450 0.8325 1.6050 0.8925 ;
        RECT 1.4400 0.4800 1.5000 0.5400 ;
        RECT 1.3350 0.3000 1.3950 0.3600 ;
        RECT 1.3350 0.6750 1.3950 0.7350 ;
        RECT 1.2300 0.4800 1.2900 0.5400 ;
        RECT 1.1250 0.1575 1.1850 0.2175 ;
        RECT 1.1250 0.8550 1.1850 0.9150 ;
        RECT 1.0200 0.4800 1.0800 0.5400 ;
        RECT 0.9150 0.3000 0.9750 0.3600 ;
        RECT 0.9150 0.6750 0.9750 0.7350 ;
        RECT 0.8100 0.4800 0.8700 0.5400 ;
        RECT 0.7050 0.1575 0.7650 0.2175 ;
        RECT 0.7050 0.8550 0.7650 0.9150 ;
        RECT 0.6000 0.4950 0.6600 0.5550 ;
        RECT 0.4950 0.3000 0.5550 0.3600 ;
        RECT 0.4950 0.6750 0.5550 0.7350 ;
        RECT 0.3900 0.4950 0.4500 0.5550 ;
        RECT 0.2850 0.1575 0.3450 0.2175 ;
        RECT 0.2850 0.8550 0.3450 0.9150 ;
        RECT 0.1875 0.4950 0.2475 0.5550 ;
        RECT 0.0750 0.3000 0.1350 0.3600 ;
        RECT 0.0750 0.7800 0.1350 0.8400 ;
        LAYER M1 ;
        RECT 2.0625 0.4500 2.6625 0.5700 ;
        RECT 2.3775 0.1800 2.4525 0.3750 ;
        RECT 2.0325 0.3000 2.3775 0.3750 ;
        RECT 1.9575 0.1500 2.0325 0.3750 ;
        RECT 1.5150 0.1500 1.9575 0.2250 ;
        RECT 1.8225 0.4650 1.9425 0.5700 ;
        RECT 0.8850 0.3000 1.8450 0.3750 ;
        RECT 1.4325 0.4500 1.8225 0.5700 ;
        RECT 0.8025 0.4500 1.3125 0.5700 ;
        RECT 0.2550 0.1500 1.2825 0.2250 ;
        RECT 0.1875 0.4650 0.6900 0.5850 ;
    END
END ND4_0001


MACRO ND4_0011
    CLASS CORE ;
    FOREIGN ND4_0011 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.1000 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 1.7325 0.6675 1.8375 0.8325 ;
        RECT 1.4175 0.6675 1.7325 0.7500 ;
        RECT 1.3125 0.6675 1.4175 0.8325 ;
        RECT 0.7875 0.6675 1.3125 0.7500 ;
        RECT 0.6825 0.6675 0.7875 0.8325 ;
        RECT 0.6000 0.6675 0.6825 0.7500 ;
        RECT 0.3675 0.6750 0.6000 0.7500 ;
        RECT 0.2550 0.3000 0.3750 0.4050 ;
        RECT 0.2625 0.6750 0.3675 0.8325 ;
        RECT 0.1125 0.6750 0.2625 0.7575 ;
        RECT 0.1125 0.3300 0.2550 0.4050 ;
        RECT 0.0375 0.3300 0.1125 0.7575 ;
        END
    END ZN
    PIN A4
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.6425 0.2625 1.7475 0.6075 ;
        RECT 1.1775 0.2625 1.6425 0.3375 ;
        VIA 1.6950 0.5250 VIA12_square ;
        END
    END A4
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.3725 0.5625 1.5000 0.6375 ;
        RECT 1.2075 0.4800 1.3725 0.6375 ;
        RECT 1.0350 0.5625 1.2075 0.6375 ;
        VIA 1.2900 0.5325 VIA12_square ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.7875 0.4125 1.0425 0.4875 ;
        RECT 0.6825 0.4125 0.7875 0.6150 ;
        RECT 0.5775 0.4125 0.6825 0.4875 ;
        VIA 0.7350 0.5325 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.4575 0.2625 0.9225 0.3375 ;
        RECT 0.3525 0.2625 0.4575 0.6075 ;
        VIA 0.4050 0.5250 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.8375 -0.0750 2.1000 0.0750 ;
        RECT 1.7325 -0.0750 1.8375 0.2250 ;
        RECT 0.0000 -0.0750 1.7325 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 2.0325 0.9750 2.1000 1.1250 ;
        RECT 1.9575 0.8025 2.0325 1.1250 ;
        RECT 1.6275 0.9750 1.9575 1.1250 ;
        RECT 1.5225 0.8325 1.6275 1.1250 ;
        RECT 1.2150 0.9750 1.5225 1.1250 ;
        RECT 1.0950 0.8325 1.2150 1.1250 ;
        RECT 1.0050 0.9750 1.0950 1.1250 ;
        RECT 0.8850 0.8325 1.0050 1.1250 ;
        RECT 0.5775 0.9750 0.8850 1.1250 ;
        RECT 0.4725 0.8325 0.5775 1.1250 ;
        RECT 0.1650 0.9750 0.4725 1.1250 ;
        RECT 0.0450 0.8325 0.1650 1.1250 ;
        RECT 0.0000 0.9750 0.0450 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.9650 0.2175 2.0250 0.2775 ;
        RECT 1.9650 0.8325 2.0250 0.8925 ;
        RECT 1.8600 0.4800 1.9200 0.5400 ;
        RECT 1.7550 0.1425 1.8150 0.2025 ;
        RECT 1.7550 0.7500 1.8150 0.8100 ;
        RECT 1.6500 0.4800 1.7100 0.5400 ;
        RECT 1.5450 0.2400 1.6050 0.3000 ;
        RECT 1.5450 0.8550 1.6050 0.9150 ;
        RECT 1.4400 0.4950 1.5000 0.5550 ;
        RECT 1.3350 0.3150 1.3950 0.3750 ;
        RECT 1.3350 0.7500 1.3950 0.8100 ;
        RECT 1.2300 0.4950 1.2900 0.5550 ;
        RECT 1.1250 0.1725 1.1850 0.2325 ;
        RECT 1.1250 0.8325 1.1850 0.8925 ;
        RECT 0.9150 0.1725 0.9750 0.2325 ;
        RECT 0.9150 0.8325 0.9750 0.8925 ;
        RECT 0.8100 0.4950 0.8700 0.5550 ;
        RECT 0.7050 0.3150 0.7650 0.3750 ;
        RECT 0.7050 0.7500 0.7650 0.8100 ;
        RECT 0.6000 0.4950 0.6600 0.5550 ;
        RECT 0.4950 0.1575 0.5550 0.2175 ;
        RECT 0.4950 0.8625 0.5550 0.9225 ;
        RECT 0.3900 0.4950 0.4500 0.5550 ;
        RECT 0.2850 0.3225 0.3450 0.3825 ;
        RECT 0.2850 0.7500 0.3450 0.8100 ;
        RECT 0.1875 0.5100 0.2475 0.5700 ;
        RECT 0.0750 0.1725 0.1350 0.2325 ;
        RECT 0.0750 0.8325 0.1350 0.8925 ;
        LAYER M1 ;
        RECT 1.9575 0.1800 2.0325 0.3750 ;
        RECT 1.6125 0.4500 1.9650 0.5700 ;
        RECT 1.6125 0.3000 1.9575 0.3750 ;
        RECT 1.5375 0.1500 1.6125 0.3750 ;
        RECT 1.2075 0.1500 1.5375 0.2250 ;
        RECT 1.4025 0.4650 1.5075 0.5925 ;
        RECT 1.3350 0.3150 1.4250 0.3900 ;
        RECT 1.1175 0.4875 1.4025 0.5925 ;
        RECT 1.2600 0.3150 1.3350 0.4125 ;
        RECT 0.8475 0.3375 1.2600 0.4125 ;
        RECT 1.1025 0.1500 1.2075 0.2550 ;
        RECT 0.8925 0.1500 0.9975 0.2550 ;
        RECT 0.7050 0.4875 0.9825 0.5850 ;
        RECT 0.1575 0.1500 0.8925 0.2250 ;
        RECT 0.7725 0.3150 0.8475 0.4125 ;
        RECT 0.6750 0.3150 0.7725 0.3900 ;
        RECT 0.6000 0.4650 0.7050 0.5850 ;
        RECT 0.1875 0.4800 0.4950 0.6000 ;
        RECT 0.0525 0.1500 0.1575 0.2550 ;
    END
END ND4_0011


MACRO ND4_0100
    CLASS CORE ;
    FOREIGN ND4_0100 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.3600 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 1.9425 0.2625 2.1000 0.3825 ;
        RECT 1.9425 0.6600 2.1000 0.7800 ;
        RECT 1.6275 0.2625 1.9425 0.7800 ;
        RECT 1.4700 0.2625 1.6275 0.3825 ;
        RECT 1.4700 0.6600 1.6275 0.7800 ;
        VIA 1.9425 0.3225 VIA12_slot ;
        VIA 1.9425 0.7200 VIA12_slot ;
        VIA 1.6275 0.3225 VIA12_slot ;
        VIA 1.6275 0.7200 VIA12_slot ;
        END
    END ZN
    PIN A4
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.7275 0.5625 1.2600 0.6375 ;
        VIA 0.9075 0.6000 VIA12_square ;
        END
    END A4
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.5175 0.2625 0.9825 0.3375 ;
        VIA 0.7275 0.3000 VIA12_square ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.4725 0.8625 0.6600 0.9375 ;
        RECT 0.3975 0.4050 0.4725 0.9375 ;
        RECT 0.1200 0.8625 0.3975 0.9375 ;
        VIA 0.4350 0.5100 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.3375 0.1125 0.6075 0.1875 ;
        RECT 0.2625 0.1125 0.3375 0.2775 ;
        RECT 0.0675 0.1125 0.2625 0.1875 ;
        VIA 0.3000 0.1950 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 3.1050 -0.0750 3.3600 0.0750 ;
        RECT 2.9850 -0.0750 3.1050 0.1875 ;
        RECT 2.6850 -0.0750 2.9850 0.0750 ;
        RECT 2.5650 -0.0750 2.6850 0.1875 ;
        RECT 2.2650 -0.0750 2.5650 0.0750 ;
        RECT 2.1450 -0.0750 2.2650 0.1875 ;
        RECT 1.8450 -0.0750 2.1450 0.0750 ;
        RECT 1.7250 -0.0750 1.8450 0.1875 ;
        RECT 1.4250 -0.0750 1.7250 0.0750 ;
        RECT 1.3050 -0.0750 1.4250 0.1875 ;
        RECT 1.0050 -0.0750 1.3050 0.0750 ;
        RECT 0.8850 -0.0750 1.0050 0.2475 ;
        RECT 0.0000 -0.0750 0.8850 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 3.0975 0.9750 3.3600 1.1250 ;
        RECT 2.9925 0.8100 3.0975 1.1250 ;
        RECT 2.6850 0.9750 2.9925 1.1250 ;
        RECT 2.5650 0.8175 2.6850 1.1250 ;
        RECT 2.2650 0.9750 2.5650 1.1250 ;
        RECT 2.1450 0.8550 2.2650 1.1250 ;
        RECT 1.8450 0.9750 2.1450 1.1250 ;
        RECT 1.7250 0.8550 1.8450 1.1250 ;
        RECT 1.4250 0.9750 1.7250 1.1250 ;
        RECT 1.3050 0.8550 1.4250 1.1250 ;
        RECT 1.0050 0.9750 1.3050 1.1250 ;
        RECT 0.8850 0.8025 1.0050 1.1250 ;
        RECT 0.5775 0.9750 0.8850 1.1250 ;
        RECT 0.4725 0.8475 0.5775 1.1250 ;
        RECT 0.1650 0.9750 0.4725 1.1250 ;
        RECT 0.0450 0.8175 0.1650 1.1250 ;
        RECT 0.0000 0.9750 0.0450 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 3.2250 0.2250 3.2850 0.2850 ;
        RECT 3.2250 0.7575 3.2850 0.8175 ;
        RECT 3.1200 0.4650 3.1800 0.5250 ;
        RECT 3.0150 0.1275 3.0750 0.1875 ;
        RECT 3.0150 0.8325 3.0750 0.8925 ;
        RECT 2.9100 0.4650 2.9700 0.5250 ;
        RECT 2.8050 0.2700 2.8650 0.3300 ;
        RECT 2.8050 0.6675 2.8650 0.7275 ;
        RECT 2.7000 0.4650 2.7600 0.5250 ;
        RECT 2.5950 0.1275 2.6550 0.1875 ;
        RECT 2.5950 0.8250 2.6550 0.8850 ;
        RECT 2.4900 0.4650 2.5500 0.5250 ;
        RECT 2.3850 0.2850 2.4450 0.3450 ;
        RECT 2.3850 0.6900 2.4450 0.7500 ;
        RECT 2.2800 0.4650 2.3400 0.5250 ;
        RECT 2.1750 0.1275 2.2350 0.1875 ;
        RECT 2.1750 0.8625 2.2350 0.9225 ;
        RECT 2.0700 0.4650 2.1300 0.5250 ;
        RECT 1.9650 0.2850 2.0250 0.3450 ;
        RECT 1.9650 0.6900 2.0250 0.7500 ;
        RECT 1.8600 0.4650 1.9200 0.5250 ;
        RECT 1.7550 0.1275 1.8150 0.1875 ;
        RECT 1.7550 0.8625 1.8150 0.9225 ;
        RECT 1.6500 0.4650 1.7100 0.5250 ;
        RECT 1.5450 0.2850 1.6050 0.3450 ;
        RECT 1.5450 0.6900 1.6050 0.7500 ;
        RECT 1.4400 0.4650 1.5000 0.5250 ;
        RECT 1.3350 0.1275 1.3950 0.1875 ;
        RECT 1.3350 0.8625 1.3950 0.9225 ;
        RECT 1.2300 0.4650 1.2900 0.5250 ;
        RECT 1.1250 0.2850 1.1850 0.3450 ;
        RECT 1.1250 0.6900 1.1850 0.7500 ;
        RECT 1.0200 0.4875 1.0800 0.5475 ;
        RECT 0.9150 0.1575 0.9750 0.2175 ;
        RECT 0.9150 0.8325 0.9750 0.8925 ;
        RECT 0.8100 0.4650 0.8700 0.5250 ;
        RECT 0.7050 0.7200 0.7650 0.7800 ;
        RECT 0.6000 0.4650 0.6600 0.5250 ;
        RECT 0.4950 0.8700 0.5550 0.9300 ;
        RECT 0.3900 0.4650 0.4500 0.5250 ;
        RECT 0.2850 0.6825 0.3450 0.7425 ;
        RECT 0.1875 0.4650 0.2475 0.5250 ;
        RECT 0.0750 0.1800 0.1350 0.2400 ;
        RECT 0.0750 0.8325 0.1350 0.8925 ;
        LAYER M1 ;
        RECT 3.2025 0.1950 3.3075 0.3375 ;
        RECT 3.2175 0.6600 3.2925 0.8700 ;
        RECT 2.8050 0.4125 3.2475 0.5325 ;
        RECT 2.6175 0.6600 3.2175 0.7350 ;
        RECT 2.6175 0.2625 3.2025 0.3375 ;
        RECT 2.7000 0.4125 2.8050 0.5625 ;
        RECT 2.5425 0.2625 2.6175 0.7350 ;
        RECT 1.1250 0.4575 2.5425 0.5325 ;
        RECT 1.1025 0.2625 2.4675 0.3825 ;
        RECT 1.1025 0.6600 2.4675 0.7800 ;
        RECT 1.0200 0.4575 1.1250 0.5775 ;
        RECT 0.8475 0.4350 0.9450 0.6825 ;
        RECT 0.7800 0.4350 0.8475 0.5550 ;
        RECT 0.6975 0.2400 0.8100 0.3600 ;
        RECT 0.6900 0.6675 0.7650 0.8325 ;
        RECT 0.5925 0.2400 0.6975 0.5550 ;
        RECT 0.1125 0.6675 0.6900 0.7425 ;
        RECT 0.3675 0.3600 0.5175 0.5925 ;
        RECT 0.2925 0.1500 0.3825 0.2475 ;
        RECT 0.2175 0.1500 0.2925 0.5550 ;
        RECT 0.1875 0.4350 0.2175 0.5550 ;
        RECT 0.1125 0.1500 0.1425 0.2700 ;
        RECT 0.0375 0.1500 0.1125 0.7425 ;
        LAYER VIA1 ;
        RECT 2.7975 0.4125 2.8725 0.4875 ;
        RECT 0.6900 0.7125 0.7650 0.7875 ;
        LAYER M2 ;
        RECT 1.9725 0.2625 2.1000 0.3825 ;
        RECT 1.9725 0.6600 2.1000 0.7800 ;
        RECT 1.4700 0.2625 1.5975 0.3825 ;
        RECT 1.4700 0.6600 1.5975 0.7800 ;
        RECT 2.3250 0.4125 3.0075 0.4875 ;
        RECT 2.2500 0.4125 2.3250 0.9375 ;
        RECT 1.0275 0.8625 2.2500 0.9375 ;
        RECT 0.9525 0.7125 1.0275 0.9375 ;
        RECT 0.6375 0.7125 0.9525 0.7875 ;
    END
END ND4_0100


MACRO ND4_0111
    CLASS CORE ;
    FOREIGN ND4_0111 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.7800 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 0.3675 0.2700 0.6825 0.8025 ;
        VIA 0.5250 0.3525 VIA12_slot ;
        VIA 0.5250 0.7200 VIA12_slot ;
        END
    END ZN
    PIN A4
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 3.1425 0.4125 3.2475 0.6225 ;
        RECT 2.6775 0.4125 3.1425 0.4875 ;
        VIA 3.1950 0.5175 VIA12_square ;
        END
    END A4
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 2.3850 0.4125 2.4900 0.6225 ;
        RECT 1.9200 0.4125 2.3850 0.4875 ;
        VIA 2.4375 0.5400 VIA12_square ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.5225 0.4125 1.6275 0.6225 ;
        RECT 1.0575 0.4125 1.5225 0.4875 ;
        VIA 1.5750 0.5400 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1725 0.4800 0.9075 0.5850 ;
        RECT 0.1425 0.4800 0.1725 0.6825 ;
        RECT 0.0675 0.3675 0.1425 0.6825 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 3.5175 -0.0750 3.7800 0.0750 ;
        RECT 3.4125 -0.0750 3.5175 0.2250 ;
        RECT 3.0975 -0.0750 3.4125 0.0750 ;
        RECT 2.9925 -0.0750 3.0975 0.2250 ;
        RECT 0.0000 -0.0750 2.9925 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 3.7125 0.9750 3.7800 1.1250 ;
        RECT 3.6375 0.8025 3.7125 1.1250 ;
        RECT 3.3075 0.9750 3.6375 1.1250 ;
        RECT 3.2025 0.8325 3.3075 1.1250 ;
        RECT 2.8875 0.9750 3.2025 1.1250 ;
        RECT 2.7825 0.8325 2.8875 1.1250 ;
        RECT 2.4675 0.9750 2.7825 1.1250 ;
        RECT 2.3625 0.8325 2.4675 1.1250 ;
        RECT 2.0550 0.9750 2.3625 1.1250 ;
        RECT 1.9350 0.8325 2.0550 1.1250 ;
        RECT 1.8450 0.9750 1.9350 1.1250 ;
        RECT 1.7250 0.8325 1.8450 1.1250 ;
        RECT 1.4175 0.9750 1.7250 1.1250 ;
        RECT 1.3125 0.8325 1.4175 1.1250 ;
        RECT 0.9975 0.9750 1.3125 1.1250 ;
        RECT 0.8925 0.8325 0.9975 1.1250 ;
        RECT 0.5775 0.9750 0.8925 1.1250 ;
        RECT 0.4725 0.8325 0.5775 1.1250 ;
        RECT 0.1425 0.9750 0.4725 1.1250 ;
        RECT 0.0675 0.8025 0.1425 1.1250 ;
        RECT 0.0000 0.9750 0.0675 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 3.6450 0.2175 3.7050 0.2775 ;
        RECT 3.6450 0.8325 3.7050 0.8925 ;
        RECT 3.5400 0.4800 3.6000 0.5400 ;
        RECT 3.4350 0.1425 3.4950 0.2025 ;
        RECT 3.4350 0.6900 3.4950 0.7500 ;
        RECT 3.3300 0.4800 3.3900 0.5400 ;
        RECT 3.2250 0.3000 3.2850 0.3600 ;
        RECT 3.2250 0.8550 3.2850 0.9150 ;
        RECT 3.1200 0.4800 3.1800 0.5400 ;
        RECT 3.0150 0.1425 3.0750 0.2025 ;
        RECT 3.0150 0.6900 3.0750 0.7500 ;
        RECT 2.9100 0.4800 2.9700 0.5400 ;
        RECT 2.8050 0.2400 2.8650 0.3000 ;
        RECT 2.8050 0.8550 2.8650 0.9150 ;
        RECT 2.7000 0.4950 2.7600 0.5550 ;
        RECT 2.5950 0.3150 2.6550 0.3750 ;
        RECT 2.5950 0.6900 2.6550 0.7500 ;
        RECT 2.4900 0.4950 2.5500 0.5550 ;
        RECT 2.3850 0.1575 2.4450 0.2175 ;
        RECT 2.3850 0.8550 2.4450 0.9150 ;
        RECT 2.2800 0.4950 2.3400 0.5550 ;
        RECT 2.1750 0.3150 2.2350 0.3750 ;
        RECT 2.1750 0.6900 2.2350 0.7500 ;
        RECT 2.0700 0.4950 2.1300 0.5550 ;
        RECT 1.9650 0.1725 2.0250 0.2325 ;
        RECT 1.9650 0.8325 2.0250 0.8925 ;
        RECT 1.7550 0.1725 1.8150 0.2325 ;
        RECT 1.7550 0.8325 1.8150 0.8925 ;
        RECT 1.6500 0.4950 1.7100 0.5550 ;
        RECT 1.5450 0.3150 1.6050 0.3750 ;
        RECT 1.5450 0.6900 1.6050 0.7500 ;
        RECT 1.4400 0.4950 1.5000 0.5550 ;
        RECT 1.3350 0.1575 1.3950 0.2175 ;
        RECT 1.3350 0.8550 1.3950 0.9150 ;
        RECT 1.2300 0.4950 1.2900 0.5550 ;
        RECT 1.1250 0.3150 1.1850 0.3750 ;
        RECT 1.1250 0.6900 1.1850 0.7500 ;
        RECT 1.0200 0.4950 1.0800 0.5550 ;
        RECT 0.9150 0.1575 0.9750 0.2175 ;
        RECT 0.9150 0.8625 0.9750 0.9225 ;
        RECT 0.8100 0.4800 0.8700 0.5400 ;
        RECT 0.7050 0.3000 0.7650 0.3600 ;
        RECT 0.7050 0.6900 0.7650 0.7500 ;
        RECT 0.6000 0.4800 0.6600 0.5400 ;
        RECT 0.4950 0.1575 0.5550 0.2175 ;
        RECT 0.4950 0.8550 0.5550 0.9150 ;
        RECT 0.3900 0.4800 0.4500 0.5400 ;
        RECT 0.2850 0.3000 0.3450 0.3600 ;
        RECT 0.2850 0.7200 0.3450 0.7800 ;
        RECT 0.1800 0.4800 0.2400 0.5400 ;
        RECT 0.0750 0.1725 0.1350 0.2325 ;
        RECT 0.0750 0.8325 0.1350 0.8925 ;
        LAYER M1 ;
        RECT 3.6375 0.1800 3.7125 0.3750 ;
        RECT 2.8725 0.3000 3.6375 0.3750 ;
        RECT 2.9025 0.4500 3.6375 0.5700 ;
        RECT 0.3675 0.6825 3.5250 0.7575 ;
        RECT 2.7975 0.1500 2.8725 0.3750 ;
        RECT 2.0475 0.1500 2.7975 0.2250 ;
        RECT 2.6625 0.4650 2.7675 0.5925 ;
        RECT 2.2125 0.3150 2.6850 0.3900 ;
        RECT 1.9575 0.4875 2.6625 0.5925 ;
        RECT 2.1375 0.3150 2.2125 0.4125 ;
        RECT 1.6425 0.3375 2.1375 0.4125 ;
        RECT 1.9425 0.1500 2.0475 0.2550 ;
        RECT 1.7325 0.1500 1.8375 0.2550 ;
        RECT 1.1250 0.4875 1.8225 0.5850 ;
        RECT 0.1575 0.1500 1.7325 0.2250 ;
        RECT 1.5675 0.3150 1.6425 0.4125 ;
        RECT 1.0950 0.3150 1.5675 0.3900 ;
        RECT 1.0200 0.4650 1.1250 0.5850 ;
        RECT 0.2175 0.3000 0.8100 0.4050 ;
        RECT 0.2625 0.6825 0.3675 0.8025 ;
        RECT 0.0525 0.1500 0.1575 0.2550 ;
    END
END ND4_0111


MACRO ND4_1000
    CLASS CORE ;
    FOREIGN ND4_1000 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.0500 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.9375 0.1500 1.0125 0.7425 ;
        RECT 0.9075 0.1500 0.9375 0.2700 ;
        RECT 0.7875 0.6675 0.9375 0.7425 ;
        RECT 0.6825 0.6675 0.7875 0.9000 ;
        RECT 0.3675 0.6675 0.6825 0.7425 ;
        RECT 0.2625 0.6675 0.3675 0.9000 ;
        END
    END ZN
    PIN A4
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1425 0.4350 0.2475 0.5550 ;
        RECT 0.0675 0.3675 0.1425 0.6825 ;
        END
    END A4
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.0675 0.2625 0.5325 0.3375 ;
        VIA 0.3225 0.3000 VIA12_square ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.6525 0.8625 0.9300 0.9375 ;
        RECT 0.5775 0.4050 0.6525 0.9375 ;
        RECT 0.3900 0.8625 0.5775 0.9375 ;
        VIA 0.6150 0.5100 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.7875 0.1125 0.9825 0.1875 ;
        RECT 0.7125 0.1125 0.7875 0.2775 ;
        RECT 0.4425 0.1125 0.7125 0.1875 ;
        VIA 0.7500 0.1950 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.1650 -0.0750 1.0500 0.0750 ;
        RECT 0.0450 -0.0750 0.1650 0.2475 ;
        RECT 0.0000 -0.0750 0.0450 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.0050 0.9750 1.0500 1.1250 ;
        RECT 0.8850 0.8175 1.0050 1.1250 ;
        RECT 0.5775 0.9750 0.8850 1.1250 ;
        RECT 0.4725 0.8475 0.5775 1.1250 ;
        RECT 0.1650 0.9750 0.4725 1.1250 ;
        RECT 0.0450 0.8025 0.1650 1.1250 ;
        RECT 0.0000 0.9750 0.0450 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 0.9150 0.1800 0.9750 0.2400 ;
        RECT 0.9150 0.8325 0.9750 0.8925 ;
        RECT 0.8025 0.4650 0.8625 0.5250 ;
        RECT 0.7050 0.8175 0.7650 0.8775 ;
        RECT 0.6000 0.4650 0.6600 0.5250 ;
        RECT 0.4950 0.8700 0.5550 0.9300 ;
        RECT 0.3900 0.4650 0.4500 0.5250 ;
        RECT 0.2850 0.8175 0.3450 0.8775 ;
        RECT 0.1800 0.4650 0.2400 0.5250 ;
        RECT 0.0750 0.1575 0.1350 0.2175 ;
        RECT 0.0750 0.8325 0.1350 0.8925 ;
        LAYER M1 ;
        RECT 0.8325 0.4350 0.8625 0.5550 ;
        RECT 0.7575 0.1500 0.8325 0.5550 ;
        RECT 0.6675 0.1500 0.7575 0.2475 ;
        RECT 0.5325 0.3600 0.6825 0.5925 ;
        RECT 0.3225 0.2400 0.4575 0.5550 ;
        RECT 0.2400 0.2400 0.3225 0.3600 ;
    END
END ND4_1000


MACRO ND4_1010
    CLASS CORE ;
    FOREIGN ND4_1010 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.0500 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.9375 0.1500 1.0125 0.7050 ;
        RECT 0.9075 0.1500 0.9375 0.2700 ;
        RECT 0.8325 0.6300 0.9375 0.7050 ;
        RECT 0.7575 0.6300 0.8325 0.7875 ;
        RECT 0.3675 0.7125 0.7575 0.7875 ;
        RECT 0.2550 0.7125 0.3675 0.8175 ;
        END
    END ZN
    PIN A4
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1425 0.4350 0.2475 0.5550 ;
        RECT 0.0675 0.3675 0.1425 0.6825 ;
        END
    END A4
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.3375 0.2175 0.4425 0.5775 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.5175 0.3600 0.6825 0.6375 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.8325 0.3450 0.8625 0.5550 ;
        RECT 0.7575 0.2175 0.8325 0.5550 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.1650 -0.0750 1.0500 0.0750 ;
        RECT 0.0450 -0.0750 0.1650 0.2475 ;
        RECT 0.0000 -0.0750 0.0450 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.0125 0.9750 1.0500 1.1250 ;
        RECT 0.9075 0.8025 1.0125 1.1250 ;
        RECT 0.5850 0.9750 0.9075 1.1250 ;
        RECT 0.4650 0.8625 0.5850 1.1250 ;
        RECT 0.1650 0.9750 0.4650 1.1250 ;
        RECT 0.0450 0.8025 0.1650 1.1250 ;
        RECT 0.0000 0.9750 0.0450 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 0.9150 0.1800 0.9750 0.2400 ;
        RECT 0.9150 0.8325 0.9750 0.8925 ;
        RECT 0.8025 0.4650 0.8625 0.5250 ;
        RECT 0.7050 0.7200 0.7650 0.7800 ;
        RECT 0.6000 0.4650 0.6600 0.5250 ;
        RECT 0.4950 0.8700 0.5550 0.9300 ;
        RECT 0.3825 0.4650 0.4425 0.5250 ;
        RECT 0.2850 0.7350 0.3450 0.7950 ;
        RECT 0.1800 0.4650 0.2400 0.5250 ;
        RECT 0.0750 0.1725 0.1350 0.2325 ;
        RECT 0.0750 0.8325 0.1350 0.8925 ;
    END
END ND4_1010


MACRO NR2_0001
    CLASS CORE ;
    FOREIGN NR2_0001 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.4700 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.2550 0.2850 1.2150 0.3750 ;
        RECT 0.1125 0.8175 0.5850 0.9000 ;
        RECT 0.1125 0.3000 0.2550 0.3750 ;
        RECT 0.0375 0.3000 0.1125 0.9000 ;
        END
    END ZN
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.3275 0.3675 1.4025 0.6825 ;
        RECT 0.7875 0.4650 1.3275 0.5700 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.5775 0.5625 0.9525 0.6375 ;
        RECT 0.4725 0.4425 0.5775 0.6375 ;
        VIA 0.5250 0.5175 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.4025 -0.0750 1.4700 0.0750 ;
        RECT 1.3275 -0.0750 1.4025 0.2475 ;
        RECT 1.0050 -0.0750 1.3275 0.0750 ;
        RECT 0.8850 -0.0750 1.0050 0.2100 ;
        RECT 0.5850 -0.0750 0.8850 0.0750 ;
        RECT 0.4650 -0.0750 0.5850 0.2100 ;
        RECT 0.1650 -0.0750 0.4650 0.0750 ;
        RECT 0.0450 -0.0750 0.1650 0.2250 ;
        RECT 0.0000 -0.0750 0.0450 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.4250 0.9750 1.4700 1.1250 ;
        RECT 1.3050 0.7950 1.4250 1.1250 ;
        RECT 0.9975 0.9750 1.3050 1.1250 ;
        RECT 0.8925 0.8175 0.9975 1.1250 ;
        RECT 0.0000 0.9750 0.8925 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.3350 0.1575 1.3950 0.2175 ;
        RECT 1.3350 0.8325 1.3950 0.8925 ;
        RECT 1.2300 0.4875 1.2900 0.5475 ;
        RECT 1.1250 0.2925 1.1850 0.3525 ;
        RECT 1.1250 0.6900 1.1850 0.7500 ;
        RECT 1.0200 0.4875 1.0800 0.5475 ;
        RECT 0.9150 0.1425 0.9750 0.2025 ;
        RECT 0.9150 0.8400 0.9750 0.9000 ;
        RECT 0.8100 0.4875 0.8700 0.5475 ;
        RECT 0.7050 0.2925 0.7650 0.3525 ;
        RECT 0.7050 0.6825 0.7650 0.7425 ;
        RECT 0.6000 0.4725 0.6600 0.5325 ;
        RECT 0.4950 0.1425 0.5550 0.2025 ;
        RECT 0.4950 0.8250 0.5550 0.8850 ;
        RECT 0.3900 0.4725 0.4500 0.5325 ;
        RECT 0.2850 0.2925 0.3450 0.3525 ;
        RECT 0.2850 0.6750 0.3450 0.7350 ;
        RECT 0.1875 0.4950 0.2475 0.5550 ;
        RECT 0.0750 0.1575 0.1350 0.2175 ;
        RECT 0.0750 0.8250 0.1350 0.8850 ;
        LAYER M1 ;
        RECT 1.1025 0.6675 1.2075 0.7725 ;
        RECT 0.2550 0.6675 1.1025 0.7425 ;
        RECT 0.2925 0.4650 0.6900 0.5700 ;
        RECT 0.1875 0.4650 0.2925 0.5850 ;
    END
END NR2_0001


MACRO NR2_0010
    CLASS CORE ;
    FOREIGN NR2_0010 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.4100 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 1.5225 0.2850 1.6800 0.4050 ;
        RECT 1.5225 0.6375 1.6800 0.7575 ;
        RECT 1.2075 0.2850 1.5225 0.7575 ;
        RECT 1.0500 0.2850 1.2075 0.4050 ;
        RECT 1.0500 0.6375 1.2075 0.7575 ;
        VIA 1.5225 0.3450 VIA12_slot ;
        VIA 1.5225 0.6975 VIA12_slot ;
        VIA 1.2075 0.3450 VIA12_slot ;
        VIA 1.2075 0.6975 VIA12_slot ;
        END
    END ZN
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 4.0725 0.4125 4.2375 0.6375 ;
        RECT 1.8300 0.4575 4.0725 0.5775 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1575 0.4650 1.7400 0.5700 ;
        RECT 0.0525 0.3675 0.1575 0.6825 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 4.3425 -0.0750 4.4100 0.0750 ;
        RECT 4.2675 -0.0750 4.3425 0.2700 ;
        RECT 3.9450 -0.0750 4.2675 0.0750 ;
        RECT 3.8250 -0.0750 3.9450 0.1875 ;
        RECT 3.5250 -0.0750 3.8250 0.0750 ;
        RECT 3.4050 -0.0750 3.5250 0.1875 ;
        RECT 3.1050 -0.0750 3.4050 0.0750 ;
        RECT 2.9850 -0.0750 3.1050 0.1875 ;
        RECT 2.6850 -0.0750 2.9850 0.0750 ;
        RECT 2.5650 -0.0750 2.6850 0.1875 ;
        RECT 2.2650 -0.0750 2.5650 0.0750 ;
        RECT 2.1450 -0.0750 2.2650 0.1875 ;
        RECT 1.8450 -0.0750 2.1450 0.0750 ;
        RECT 1.7250 -0.0750 1.8450 0.1875 ;
        RECT 1.4250 -0.0750 1.7250 0.0750 ;
        RECT 1.3050 -0.0750 1.4250 0.1875 ;
        RECT 1.0050 -0.0750 1.3050 0.0750 ;
        RECT 0.8850 -0.0750 1.0050 0.1875 ;
        RECT 0.5850 -0.0750 0.8850 0.0750 ;
        RECT 0.4650 -0.0750 0.5850 0.1875 ;
        RECT 0.1575 -0.0750 0.4650 0.0750 ;
        RECT 0.0525 -0.0750 0.1575 0.2625 ;
        RECT 0.0000 -0.0750 0.0525 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 4.1550 0.9750 4.4100 1.1250 ;
        RECT 4.0350 0.8625 4.1550 1.1250 ;
        RECT 3.7350 0.9750 4.0350 1.1250 ;
        RECT 3.6150 0.8625 3.7350 1.1250 ;
        RECT 3.3150 0.9750 3.6150 1.1250 ;
        RECT 3.1950 0.8625 3.3150 1.1250 ;
        RECT 2.8950 0.9750 3.1950 1.1250 ;
        RECT 2.7750 0.8625 2.8950 1.1250 ;
        RECT 2.4750 0.9750 2.7750 1.1250 ;
        RECT 2.3550 0.8625 2.4750 1.1250 ;
        RECT 2.0550 0.9750 2.3550 1.1250 ;
        RECT 1.9350 0.8625 2.0550 1.1250 ;
        RECT 0.0000 0.9750 1.9350 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 4.2750 0.1575 4.3350 0.2175 ;
        RECT 4.2750 0.7800 4.3350 0.8400 ;
        RECT 4.1700 0.4875 4.2300 0.5475 ;
        RECT 4.0650 0.1725 4.1250 0.2325 ;
        RECT 4.0650 0.8625 4.1250 0.9225 ;
        RECT 3.9600 0.4875 4.0200 0.5475 ;
        RECT 3.8550 0.1275 3.9150 0.1875 ;
        RECT 3.8550 0.7200 3.9150 0.7800 ;
        RECT 3.7500 0.4875 3.8100 0.5475 ;
        RECT 3.6450 0.1725 3.7050 0.2325 ;
        RECT 3.6450 0.8625 3.7050 0.9225 ;
        RECT 3.5400 0.4875 3.6000 0.5475 ;
        RECT 3.4350 0.1275 3.4950 0.1875 ;
        RECT 3.4350 0.7200 3.4950 0.7800 ;
        RECT 3.3300 0.4875 3.3900 0.5475 ;
        RECT 3.2250 0.1725 3.2850 0.2325 ;
        RECT 3.2250 0.8625 3.2850 0.9225 ;
        RECT 3.1200 0.4875 3.1800 0.5475 ;
        RECT 3.0150 0.1275 3.0750 0.1875 ;
        RECT 3.0150 0.7200 3.0750 0.7800 ;
        RECT 2.9100 0.4875 2.9700 0.5475 ;
        RECT 2.8050 0.1725 2.8650 0.2325 ;
        RECT 2.8050 0.8625 2.8650 0.9225 ;
        RECT 2.7000 0.4875 2.7600 0.5475 ;
        RECT 2.5950 0.1275 2.6550 0.1875 ;
        RECT 2.5950 0.7200 2.6550 0.7800 ;
        RECT 2.4900 0.4875 2.5500 0.5475 ;
        RECT 2.3850 0.2925 2.4450 0.3525 ;
        RECT 2.3850 0.8625 2.4450 0.9225 ;
        RECT 2.2800 0.4875 2.3400 0.5475 ;
        RECT 2.1750 0.1275 2.2350 0.1875 ;
        RECT 2.1750 0.7200 2.2350 0.7800 ;
        RECT 2.0700 0.4875 2.1300 0.5475 ;
        RECT 1.9650 0.2925 2.0250 0.3525 ;
        RECT 1.9650 0.8625 2.0250 0.9225 ;
        RECT 1.8600 0.4875 1.9200 0.5475 ;
        RECT 1.7550 0.1275 1.8150 0.1875 ;
        RECT 1.7550 0.8325 1.8150 0.8925 ;
        RECT 1.6500 0.4875 1.7100 0.5475 ;
        RECT 1.5450 0.2925 1.6050 0.3525 ;
        RECT 1.5450 0.6750 1.6050 0.7350 ;
        RECT 1.4400 0.4875 1.5000 0.5475 ;
        RECT 1.3350 0.1275 1.3950 0.1875 ;
        RECT 1.3350 0.8325 1.3950 0.8925 ;
        RECT 1.2300 0.4875 1.2900 0.5475 ;
        RECT 1.1250 0.2925 1.1850 0.3525 ;
        RECT 1.1250 0.6750 1.1850 0.7350 ;
        RECT 1.0200 0.4875 1.0800 0.5475 ;
        RECT 0.9150 0.1275 0.9750 0.1875 ;
        RECT 0.9150 0.8325 0.9750 0.8925 ;
        RECT 0.8100 0.4875 0.8700 0.5475 ;
        RECT 0.7050 0.2925 0.7650 0.3525 ;
        RECT 0.7050 0.6750 0.7650 0.7350 ;
        RECT 0.6000 0.4875 0.6600 0.5475 ;
        RECT 0.4950 0.1275 0.5550 0.1875 ;
        RECT 0.4950 0.8325 0.5550 0.8925 ;
        RECT 0.3900 0.4875 0.4500 0.5475 ;
        RECT 0.2850 0.2925 0.3450 0.3525 ;
        RECT 0.2850 0.6750 0.3450 0.7350 ;
        RECT 0.1800 0.4875 0.2400 0.5475 ;
        RECT 0.0750 0.1725 0.1350 0.2325 ;
        RECT 0.0750 0.8100 0.1350 0.8700 ;
        LAYER M1 ;
        RECT 4.2675 0.7125 4.3425 0.8700 ;
        RECT 1.8525 0.7125 4.2675 0.7875 ;
        RECT 4.0425 0.1500 4.1475 0.3375 ;
        RECT 3.9975 0.2625 4.0425 0.3375 ;
        RECT 3.7275 0.2625 3.9975 0.3825 ;
        RECT 3.6225 0.1500 3.7275 0.3825 ;
        RECT 3.3075 0.2625 3.6225 0.3825 ;
        RECT 3.2025 0.1500 3.3075 0.3825 ;
        RECT 2.8875 0.2625 3.2025 0.3825 ;
        RECT 2.7825 0.1500 2.8875 0.3825 ;
        RECT 0.2775 0.2625 2.7825 0.3825 ;
        RECT 1.7775 0.7125 1.8525 0.9000 ;
        RECT 0.1575 0.8250 1.7775 0.9000 ;
        RECT 0.2550 0.6450 1.7025 0.7500 ;
        RECT 0.0525 0.7800 0.1575 0.9000 ;
        LAYER M2 ;
        RECT 1.5525 0.2850 1.6800 0.4050 ;
        RECT 1.5525 0.6375 1.6800 0.7575 ;
        RECT 1.0500 0.2850 1.1775 0.4050 ;
        RECT 1.0500 0.6375 1.1775 0.7575 ;
    END
END NR2_0010


MACRO NR2_0011
    CLASS CORE ;
    FOREIGN NR2_0011 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.0500 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.6975 0.2175 0.7725 0.3825 ;
        RECT 0.6675 0.3000 0.6975 0.3825 ;
        RECT 0.1125 0.3000 0.6675 0.3750 ;
        RECT 0.1125 0.6450 0.3750 0.7200 ;
        RECT 0.0375 0.3000 0.1125 0.7200 ;
        END
    END ZN
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.9075 0.3675 1.0125 0.6375 ;
        RECT 0.6825 0.4725 0.9075 0.6375 ;
        RECT 0.5700 0.4725 0.6825 0.5775 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.4650 0.7125 0.7725 0.7875 ;
        RECT 0.3600 0.4425 0.4650 0.7875 ;
        RECT 0.3075 0.7125 0.3600 0.7875 ;
        VIA 0.4125 0.5175 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.9825 -0.0750 1.0500 0.0750 ;
        RECT 0.9075 -0.0750 0.9825 0.2475 ;
        RECT 0.5850 -0.0750 0.9075 0.0750 ;
        RECT 0.4650 -0.0750 0.5850 0.2175 ;
        RECT 0.1650 -0.0750 0.4650 0.0750 ;
        RECT 0.0450 -0.0750 0.1650 0.2250 ;
        RECT 0.0000 -0.0750 0.0450 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.7950 0.9750 1.0500 1.1250 ;
        RECT 0.6750 0.8625 0.7950 1.1250 ;
        RECT 0.0000 0.9750 0.6750 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 0.9150 0.1575 0.9750 0.2175 ;
        RECT 0.9150 0.7800 0.9750 0.8400 ;
        RECT 0.8100 0.4800 0.8700 0.5400 ;
        RECT 0.7050 0.2700 0.7650 0.3300 ;
        RECT 0.7050 0.8625 0.7650 0.9225 ;
        RECT 0.6000 0.4800 0.6600 0.5400 ;
        RECT 0.4950 0.1500 0.5550 0.2100 ;
        RECT 0.4950 0.8325 0.5550 0.8925 ;
        RECT 0.3900 0.4800 0.4500 0.5400 ;
        RECT 0.2850 0.3000 0.3450 0.3600 ;
        RECT 0.2850 0.6600 0.3450 0.7200 ;
        RECT 0.1875 0.4800 0.2475 0.5400 ;
        RECT 0.0750 0.1575 0.1350 0.2175 ;
        RECT 0.0750 0.8175 0.1350 0.8775 ;
        LAYER M1 ;
        RECT 0.9075 0.7125 0.9825 0.8700 ;
        RECT 0.6000 0.7125 0.9075 0.7875 ;
        RECT 0.5250 0.7125 0.6000 0.9000 ;
        RECT 0.1650 0.8250 0.5250 0.9000 ;
        RECT 0.1875 0.4500 0.4950 0.5700 ;
        RECT 0.0450 0.7950 0.1650 0.9000 ;
    END
END NR2_0011


MACRO NR2_0100
    CLASS CORE ;
    FOREIGN NR2_0100 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.5700 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 1.1025 0.2700 1.2600 0.3900 ;
        RECT 1.1025 0.6300 1.2600 0.7500 ;
        RECT 0.7875 0.2700 1.1025 0.7500 ;
        RECT 0.6300 0.2700 0.7875 0.3900 ;
        RECT 0.6300 0.6300 0.7875 0.7500 ;
        VIA 1.1025 0.3300 VIA12_slot ;
        VIA 1.1025 0.6900 VIA12_slot ;
        VIA 0.7875 0.3300 VIA12_slot ;
        VIA 0.7875 0.6900 VIA12_slot ;
        END
    END ZN
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 2.2575 0.4125 2.8350 0.4875 ;
        RECT 2.1525 0.4125 2.2575 0.6075 ;
        VIA 2.2050 0.5325 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1425 0.4725 1.7400 0.5475 ;
        RECT 0.0675 0.3675 0.1425 0.6825 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 3.5175 -0.0750 3.5700 0.0750 ;
        RECT 3.4125 -0.0750 3.5175 0.2625 ;
        RECT 3.1050 -0.0750 3.4125 0.0750 ;
        RECT 2.9850 -0.0750 3.1050 0.1950 ;
        RECT 2.6850 -0.0750 2.9850 0.0750 ;
        RECT 2.5650 -0.0750 2.6850 0.1950 ;
        RECT 2.2650 -0.0750 2.5650 0.0750 ;
        RECT 2.1450 -0.0750 2.2650 0.1950 ;
        RECT 1.8450 -0.0750 2.1450 0.0750 ;
        RECT 1.7250 -0.0750 1.8450 0.1950 ;
        RECT 1.4250 -0.0750 1.7250 0.0750 ;
        RECT 1.3050 -0.0750 1.4250 0.1950 ;
        RECT 1.0050 -0.0750 1.3050 0.0750 ;
        RECT 0.8850 -0.0750 1.0050 0.1950 ;
        RECT 0.5850 -0.0750 0.8850 0.0750 ;
        RECT 0.4650 -0.0750 0.5850 0.1950 ;
        RECT 0.1425 -0.0750 0.4650 0.0750 ;
        RECT 0.0675 -0.0750 0.1425 0.2625 ;
        RECT 0.0000 -0.0750 0.0675 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 3.3150 0.9750 3.5700 1.1250 ;
        RECT 3.1950 0.8250 3.3150 1.1250 ;
        RECT 2.8950 0.9750 3.1950 1.1250 ;
        RECT 2.7750 0.8250 2.8950 1.1250 ;
        RECT 2.4750 0.9750 2.7750 1.1250 ;
        RECT 2.3550 0.8250 2.4750 1.1250 ;
        RECT 2.0550 0.9750 2.3550 1.1250 ;
        RECT 1.9350 0.8250 2.0550 1.1250 ;
        RECT 0.0000 0.9750 1.9350 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 3.4350 0.1725 3.4950 0.2325 ;
        RECT 3.4350 0.6975 3.4950 0.7575 ;
        RECT 3.3300 0.4950 3.3900 0.5550 ;
        RECT 3.2250 0.3000 3.2850 0.3600 ;
        RECT 3.2250 0.8325 3.2850 0.8925 ;
        RECT 3.1200 0.4950 3.1800 0.5550 ;
        RECT 3.0150 0.1350 3.0750 0.1950 ;
        RECT 3.0150 0.6825 3.0750 0.7425 ;
        RECT 2.9100 0.4950 2.9700 0.5550 ;
        RECT 2.8050 0.3000 2.8650 0.3600 ;
        RECT 2.8050 0.8325 2.8650 0.8925 ;
        RECT 2.7000 0.4950 2.7600 0.5550 ;
        RECT 2.5950 0.1350 2.6550 0.1950 ;
        RECT 2.5950 0.6825 2.6550 0.7425 ;
        RECT 2.4900 0.4950 2.5500 0.5550 ;
        RECT 2.3850 0.3000 2.4450 0.3600 ;
        RECT 2.3850 0.8325 2.4450 0.8925 ;
        RECT 2.2800 0.4950 2.3400 0.5550 ;
        RECT 2.1750 0.1350 2.2350 0.1950 ;
        RECT 2.1750 0.6825 2.2350 0.7425 ;
        RECT 2.0700 0.4950 2.1300 0.5550 ;
        RECT 1.9650 0.3000 2.0250 0.3600 ;
        RECT 1.9650 0.8325 2.0250 0.8925 ;
        RECT 1.8600 0.4950 1.9200 0.5550 ;
        RECT 1.7550 0.1350 1.8150 0.1950 ;
        RECT 1.7550 0.7650 1.8150 0.8250 ;
        RECT 1.6500 0.4800 1.7100 0.5400 ;
        RECT 1.5450 0.3000 1.6050 0.3600 ;
        RECT 1.5450 0.6600 1.6050 0.7200 ;
        RECT 1.4400 0.4800 1.5000 0.5400 ;
        RECT 1.3350 0.1350 1.3950 0.1950 ;
        RECT 1.3350 0.8325 1.3950 0.8925 ;
        RECT 1.2300 0.4800 1.2900 0.5400 ;
        RECT 1.1250 0.3000 1.1850 0.3600 ;
        RECT 1.1250 0.6600 1.1850 0.7200 ;
        RECT 1.0200 0.4800 1.0800 0.5400 ;
        RECT 0.9150 0.1350 0.9750 0.1950 ;
        RECT 0.9150 0.8325 0.9750 0.8925 ;
        RECT 0.8100 0.4800 0.8700 0.5400 ;
        RECT 0.7050 0.3000 0.7650 0.3600 ;
        RECT 0.7050 0.6600 0.7650 0.7200 ;
        RECT 0.6000 0.4800 0.6600 0.5400 ;
        RECT 0.4950 0.1350 0.5550 0.1950 ;
        RECT 0.4950 0.8325 0.5550 0.8925 ;
        RECT 0.3900 0.4800 0.4500 0.5400 ;
        RECT 0.2850 0.3000 0.3450 0.3600 ;
        RECT 0.2850 0.6600 0.3450 0.7200 ;
        RECT 0.1800 0.4800 0.2400 0.5400 ;
        RECT 0.0750 0.1725 0.1350 0.2325 ;
        RECT 0.0750 0.8025 0.1350 0.8625 ;
        LAYER M1 ;
        RECT 3.4125 0.6750 3.5175 0.7800 ;
        RECT 1.8525 0.4650 3.4275 0.5850 ;
        RECT 1.8225 0.6750 3.4125 0.7500 ;
        RECT 0.2550 0.2700 3.3150 0.3900 ;
        RECT 1.7475 0.6750 1.8225 0.9000 ;
        RECT 0.1575 0.8250 1.7475 0.9000 ;
        RECT 0.2550 0.6300 1.6275 0.7500 ;
        RECT 0.0525 0.7800 0.1575 0.9000 ;
        LAYER M2 ;
        RECT 1.1325 0.2700 1.2600 0.3900 ;
        RECT 1.1325 0.6300 1.2600 0.7500 ;
        RECT 0.6300 0.2700 0.7575 0.3900 ;
        RECT 0.6300 0.6300 0.7575 0.7500 ;
    END
END NR2_0100


MACRO NR2_0101
    CLASS CORE ;
    FOREIGN NR2_0101 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.2500 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 1.9425 0.2700 2.1000 0.3900 ;
        RECT 1.9425 0.6300 2.1000 0.7500 ;
        RECT 1.6275 0.2700 1.9425 0.7500 ;
        RECT 1.4700 0.2700 1.6275 0.3900 ;
        RECT 1.4700 0.6300 1.6275 0.7500 ;
        VIA 1.9425 0.3300 VIA12_slot ;
        VIA 1.9425 0.6900 VIA12_slot ;
        VIA 1.6275 0.3300 VIA12_slot ;
        VIA 1.6275 0.6900 VIA12_slot ;
        END
    END ZN
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 3.0975 0.4125 3.6750 0.4875 ;
        RECT 2.9925 0.4125 3.0975 0.6075 ;
        VIA 3.0450 0.5325 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1425 0.4725 2.5800 0.5475 ;
        RECT 0.0675 0.3675 0.1425 0.6825 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 5.1975 -0.0750 5.2500 0.0750 ;
        RECT 5.0925 -0.0750 5.1975 0.2625 ;
        RECT 4.7850 -0.0750 5.0925 0.0750 ;
        RECT 4.6650 -0.0750 4.7850 0.1950 ;
        RECT 4.3650 -0.0750 4.6650 0.0750 ;
        RECT 4.2450 -0.0750 4.3650 0.1950 ;
        RECT 3.9450 -0.0750 4.2450 0.0750 ;
        RECT 3.8250 -0.0750 3.9450 0.1950 ;
        RECT 3.5250 -0.0750 3.8250 0.0750 ;
        RECT 3.4050 -0.0750 3.5250 0.1950 ;
        RECT 3.1050 -0.0750 3.4050 0.0750 ;
        RECT 2.9850 -0.0750 3.1050 0.1950 ;
        RECT 2.6850 -0.0750 2.9850 0.0750 ;
        RECT 2.5650 -0.0750 2.6850 0.1950 ;
        RECT 2.2650 -0.0750 2.5650 0.0750 ;
        RECT 2.1450 -0.0750 2.2650 0.1950 ;
        RECT 1.8450 -0.0750 2.1450 0.0750 ;
        RECT 1.7250 -0.0750 1.8450 0.1950 ;
        RECT 1.4250 -0.0750 1.7250 0.0750 ;
        RECT 1.3050 -0.0750 1.4250 0.1950 ;
        RECT 1.0050 -0.0750 1.3050 0.0750 ;
        RECT 0.8850 -0.0750 1.0050 0.1950 ;
        RECT 0.5850 -0.0750 0.8850 0.0750 ;
        RECT 0.4650 -0.0750 0.5850 0.1950 ;
        RECT 0.1425 -0.0750 0.4650 0.0750 ;
        RECT 0.0675 -0.0750 0.1425 0.2625 ;
        RECT 0.0000 -0.0750 0.0675 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 4.9950 0.9750 5.2500 1.1250 ;
        RECT 4.8750 0.8250 4.9950 1.1250 ;
        RECT 4.5750 0.9750 4.8750 1.1250 ;
        RECT 4.4550 0.8250 4.5750 1.1250 ;
        RECT 4.1550 0.9750 4.4550 1.1250 ;
        RECT 4.0350 0.8250 4.1550 1.1250 ;
        RECT 3.7350 0.9750 4.0350 1.1250 ;
        RECT 3.6150 0.8250 3.7350 1.1250 ;
        RECT 3.3150 0.9750 3.6150 1.1250 ;
        RECT 3.1950 0.8250 3.3150 1.1250 ;
        RECT 2.8950 0.9750 3.1950 1.1250 ;
        RECT 2.7750 0.8250 2.8950 1.1250 ;
        RECT 0.0000 0.9750 2.7750 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 5.1150 0.1725 5.1750 0.2325 ;
        RECT 5.1150 0.6975 5.1750 0.7575 ;
        RECT 5.0100 0.4950 5.0700 0.5550 ;
        RECT 4.9050 0.3000 4.9650 0.3600 ;
        RECT 4.9050 0.8325 4.9650 0.8925 ;
        RECT 4.8000 0.4950 4.8600 0.5550 ;
        RECT 4.6950 0.1350 4.7550 0.1950 ;
        RECT 4.6950 0.6825 4.7550 0.7425 ;
        RECT 4.5900 0.4950 4.6500 0.5550 ;
        RECT 4.4850 0.3000 4.5450 0.3600 ;
        RECT 4.4850 0.8325 4.5450 0.8925 ;
        RECT 4.3800 0.4950 4.4400 0.5550 ;
        RECT 4.2750 0.1350 4.3350 0.1950 ;
        RECT 4.2750 0.6825 4.3350 0.7425 ;
        RECT 4.1700 0.4950 4.2300 0.5550 ;
        RECT 4.0650 0.3000 4.1250 0.3600 ;
        RECT 4.0650 0.8325 4.1250 0.8925 ;
        RECT 3.9600 0.4950 4.0200 0.5550 ;
        RECT 3.8550 0.1350 3.9150 0.1950 ;
        RECT 3.8550 0.6825 3.9150 0.7425 ;
        RECT 3.7500 0.4950 3.8100 0.5550 ;
        RECT 3.6450 0.3000 3.7050 0.3600 ;
        RECT 3.6450 0.8325 3.7050 0.8925 ;
        RECT 3.5400 0.4950 3.6000 0.5550 ;
        RECT 3.4350 0.1350 3.4950 0.1950 ;
        RECT 3.4350 0.6825 3.4950 0.7425 ;
        RECT 3.3300 0.4950 3.3900 0.5550 ;
        RECT 3.2250 0.3000 3.2850 0.3600 ;
        RECT 3.2250 0.8325 3.2850 0.8925 ;
        RECT 3.1200 0.4950 3.1800 0.5550 ;
        RECT 3.0150 0.1350 3.0750 0.1950 ;
        RECT 3.0150 0.6825 3.0750 0.7425 ;
        RECT 2.9100 0.4950 2.9700 0.5550 ;
        RECT 2.8050 0.3000 2.8650 0.3600 ;
        RECT 2.8050 0.8325 2.8650 0.8925 ;
        RECT 2.7000 0.4950 2.7600 0.5550 ;
        RECT 2.5950 0.1350 2.6550 0.1950 ;
        RECT 2.5950 0.7650 2.6550 0.8250 ;
        RECT 2.4900 0.4800 2.5500 0.5400 ;
        RECT 2.3850 0.3000 2.4450 0.3600 ;
        RECT 2.3850 0.6600 2.4450 0.7200 ;
        RECT 2.2800 0.4800 2.3400 0.5400 ;
        RECT 2.1750 0.1350 2.2350 0.1950 ;
        RECT 2.1750 0.8325 2.2350 0.8925 ;
        RECT 2.0700 0.4800 2.1300 0.5400 ;
        RECT 1.9650 0.3000 2.0250 0.3600 ;
        RECT 1.9650 0.6600 2.0250 0.7200 ;
        RECT 1.8600 0.4800 1.9200 0.5400 ;
        RECT 1.7550 0.1350 1.8150 0.1950 ;
        RECT 1.7550 0.8325 1.8150 0.8925 ;
        RECT 1.6500 0.4800 1.7100 0.5400 ;
        RECT 1.5450 0.3000 1.6050 0.3600 ;
        RECT 1.5450 0.6600 1.6050 0.7200 ;
        RECT 1.4400 0.4800 1.5000 0.5400 ;
        RECT 1.3350 0.1350 1.3950 0.1950 ;
        RECT 1.3350 0.8325 1.3950 0.8925 ;
        RECT 1.2300 0.4800 1.2900 0.5400 ;
        RECT 1.1250 0.3000 1.1850 0.3600 ;
        RECT 1.1250 0.6600 1.1850 0.7200 ;
        RECT 1.0200 0.4800 1.0800 0.5400 ;
        RECT 0.9150 0.1350 0.9750 0.1950 ;
        RECT 0.9150 0.8325 0.9750 0.8925 ;
        RECT 0.8100 0.4800 0.8700 0.5400 ;
        RECT 0.7050 0.3000 0.7650 0.3600 ;
        RECT 0.7050 0.6600 0.7650 0.7200 ;
        RECT 0.6000 0.4800 0.6600 0.5400 ;
        RECT 0.4950 0.1350 0.5550 0.1950 ;
        RECT 0.4950 0.8325 0.5550 0.8925 ;
        RECT 0.3900 0.4800 0.4500 0.5400 ;
        RECT 0.2850 0.3000 0.3450 0.3600 ;
        RECT 0.2850 0.6600 0.3450 0.7200 ;
        RECT 0.1800 0.4800 0.2400 0.5400 ;
        RECT 0.0750 0.1725 0.1350 0.2325 ;
        RECT 0.0750 0.8025 0.1350 0.8625 ;
        LAYER M1 ;
        RECT 5.0925 0.6750 5.1975 0.7800 ;
        RECT 2.6925 0.4650 5.1075 0.5850 ;
        RECT 2.6625 0.6750 5.0925 0.7500 ;
        RECT 0.2550 0.2700 4.9950 0.3900 ;
        RECT 2.5875 0.6750 2.6625 0.9000 ;
        RECT 0.1575 0.8250 2.5875 0.9000 ;
        RECT 0.2550 0.6300 2.4675 0.7500 ;
        RECT 0.0525 0.7800 0.1575 0.9000 ;
        LAYER M2 ;
        RECT 1.9725 0.2700 2.1000 0.3900 ;
        RECT 1.9725 0.6300 2.1000 0.7500 ;
        RECT 1.4700 0.2700 1.5975 0.3900 ;
        RECT 1.4700 0.6300 1.5975 0.7500 ;
    END
END NR2_0101


MACRO NR2_0111
    CLASS CORE ;
    FOREIGN NR2_0111 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.8900 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 0.3675 0.2625 0.6825 0.7575 ;
        VIA 0.5250 0.3225 VIA12_slot ;
        VIA 0.5250 0.6975 VIA12_slot ;
        END
    END ZN
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.7475 0.3675 1.8225 0.6375 ;
        RECT 0.9975 0.4875 1.7475 0.6375 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1575 0.4500 0.9000 0.5550 ;
        RECT 0.0525 0.3675 0.1575 0.6825 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.8375 -0.0750 1.8900 0.0750 ;
        RECT 1.7325 -0.0750 1.8375 0.2625 ;
        RECT 1.4250 -0.0750 1.7325 0.0750 ;
        RECT 1.3050 -0.0750 1.4250 0.1950 ;
        RECT 1.0050 -0.0750 1.3050 0.0750 ;
        RECT 0.8850 -0.0750 1.0050 0.1950 ;
        RECT 0.5850 -0.0750 0.8850 0.0750 ;
        RECT 0.4650 -0.0750 0.5850 0.1950 ;
        RECT 0.1500 -0.0750 0.4650 0.0750 ;
        RECT 0.0450 -0.0750 0.1500 0.2925 ;
        RECT 0.0000 -0.0750 0.0450 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.6350 0.9750 1.8900 1.1250 ;
        RECT 1.5150 0.8625 1.6350 1.1250 ;
        RECT 1.2150 0.9750 1.5150 1.1250 ;
        RECT 1.0950 0.8625 1.2150 1.1250 ;
        RECT 0.0000 0.9750 1.0950 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.7550 0.1725 1.8150 0.2325 ;
        RECT 1.7550 0.7425 1.8150 0.8025 ;
        RECT 1.6500 0.4950 1.7100 0.5550 ;
        RECT 1.5450 0.2625 1.6050 0.3225 ;
        RECT 1.5450 0.8625 1.6050 0.9225 ;
        RECT 1.4400 0.4950 1.5000 0.5550 ;
        RECT 1.3350 0.1275 1.3950 0.1875 ;
        RECT 1.3350 0.7200 1.3950 0.7800 ;
        RECT 1.2300 0.4950 1.2900 0.5550 ;
        RECT 1.1250 0.2775 1.1850 0.3375 ;
        RECT 1.1250 0.8625 1.1850 0.9225 ;
        RECT 1.0275 0.4950 1.0875 0.5550 ;
        RECT 0.9150 0.1275 0.9750 0.1875 ;
        RECT 0.9150 0.8325 0.9750 0.8925 ;
        RECT 0.8100 0.4800 0.8700 0.5400 ;
        RECT 0.7050 0.2775 0.7650 0.3375 ;
        RECT 0.7050 0.6675 0.7650 0.7275 ;
        RECT 0.6000 0.4800 0.6600 0.5400 ;
        RECT 0.4950 0.1275 0.5550 0.1875 ;
        RECT 0.4950 0.8325 0.5550 0.8925 ;
        RECT 0.3900 0.4800 0.4500 0.5400 ;
        RECT 0.2850 0.2775 0.3450 0.3375 ;
        RECT 0.2850 0.6675 0.3450 0.7275 ;
        RECT 0.1800 0.4800 0.2400 0.5400 ;
        RECT 0.0750 0.2025 0.1350 0.2625 ;
        RECT 0.0750 0.8025 0.1350 0.8625 ;
        LAYER M1 ;
        RECT 1.7400 0.7125 1.8300 0.8325 ;
        RECT 1.0200 0.7125 1.7400 0.7875 ;
        RECT 1.5225 0.2400 1.6275 0.3750 ;
        RECT 0.2550 0.2700 1.5225 0.3750 ;
        RECT 0.9450 0.7125 1.0200 0.9000 ;
        RECT 0.1575 0.8250 0.9450 0.9000 ;
        RECT 0.2625 0.6450 0.8700 0.7500 ;
        RECT 0.0525 0.7725 0.1575 0.9000 ;
    END
END NR2_0111


MACRO NR2_1000
    CLASS CORE ;
    FOREIGN NR2_1000 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.6300 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.5175 0.3000 0.5925 0.9000 ;
        RECT 0.3675 0.3000 0.5175 0.3750 ;
        RECT 0.4725 0.6675 0.5175 0.9000 ;
        RECT 0.2625 0.1500 0.3675 0.3750 ;
        END
    END ZN
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1425 0.4500 0.2325 0.6000 ;
        RECT 0.0675 0.3675 0.1425 0.6825 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.3825 0.4500 0.4425 0.5925 ;
        RECT 0.3075 0.4500 0.3825 0.8325 ;
        RECT 0.2775 0.6675 0.3075 0.8325 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.5925 -0.0750 0.6300 0.0750 ;
        RECT 0.4500 -0.0750 0.5925 0.2250 ;
        RECT 0.1425 -0.0750 0.4500 0.0750 ;
        RECT 0.0675 -0.0750 0.1425 0.2475 ;
        RECT 0.0000 -0.0750 0.0675 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.1425 0.9750 0.6300 1.1250 ;
        RECT 0.0675 0.8025 0.1425 1.1250 ;
        RECT 0.0000 0.9750 0.0675 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 0.4950 0.1575 0.5550 0.2175 ;
        RECT 0.4950 0.8175 0.5550 0.8775 ;
        RECT 0.3825 0.4950 0.4425 0.5550 ;
        RECT 0.2850 0.1725 0.3450 0.2325 ;
        RECT 0.1725 0.4950 0.2325 0.5550 ;
        RECT 0.0750 0.1575 0.1350 0.2175 ;
        RECT 0.0750 0.8325 0.1350 0.8925 ;
    END
END NR2_1000


MACRO NR2_1010
    CLASS CORE ;
    FOREIGN NR2_1010 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.6300 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.5175 0.3000 0.5925 0.8325 ;
        RECT 0.3525 0.3000 0.5175 0.3750 ;
        RECT 0.4875 0.6675 0.5175 0.8325 ;
        RECT 0.2775 0.2175 0.3525 0.3750 ;
        END
    END ZN
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1425 0.4500 0.2325 0.6000 ;
        RECT 0.0675 0.3675 0.1425 0.6825 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.3825 0.4500 0.4425 0.6000 ;
        RECT 0.3075 0.4500 0.3825 0.8325 ;
        RECT 0.2775 0.6675 0.3075 0.8325 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.5925 -0.0750 0.6300 0.0750 ;
        RECT 0.4500 -0.0750 0.5925 0.2250 ;
        RECT 0.1425 -0.0750 0.4500 0.0750 ;
        RECT 0.0675 -0.0750 0.1425 0.2475 ;
        RECT 0.0000 -0.0750 0.0675 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.1425 0.9750 0.6300 1.1250 ;
        RECT 0.0675 0.8025 0.1425 1.1250 ;
        RECT 0.0000 0.9750 0.0675 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 0.4950 0.1575 0.5550 0.2175 ;
        RECT 0.4950 0.7200 0.5550 0.7800 ;
        RECT 0.3825 0.4950 0.4425 0.5550 ;
        RECT 0.2850 0.2625 0.3450 0.3225 ;
        RECT 0.1725 0.4950 0.2325 0.5550 ;
        RECT 0.0750 0.1575 0.1350 0.2175 ;
        RECT 0.0750 0.8325 0.1350 0.8925 ;
    END
END NR2_1010


MACRO NR2_1100
    CLASS CORE ;
    FOREIGN NR2_1100 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.9300 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 2.7825 0.2700 2.9400 0.3900 ;
        RECT 2.7825 0.6300 2.9400 0.7500 ;
        RECT 2.4675 0.2700 2.7825 0.7500 ;
        RECT 2.3100 0.2700 2.4675 0.3900 ;
        RECT 2.3100 0.6300 2.4675 0.7500 ;
        VIA 2.7825 0.3300 VIA12_slot ;
        VIA 2.7825 0.6900 VIA12_slot ;
        VIA 2.4675 0.3300 VIA12_slot ;
        VIA 2.4675 0.6900 VIA12_slot ;
        END
    END ZN
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 4.7325 0.4125 5.3100 0.4875 ;
        RECT 4.6275 0.4125 4.7325 0.6075 ;
        VIA 4.6800 0.5325 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1425 0.4725 3.4200 0.5475 ;
        RECT 0.0675 0.3675 0.1425 0.6825 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 6.8775 -0.0750 6.9300 0.0750 ;
        RECT 6.7725 -0.0750 6.8775 0.2625 ;
        RECT 6.4650 -0.0750 6.7725 0.0750 ;
        RECT 6.3450 -0.0750 6.4650 0.1950 ;
        RECT 6.0450 -0.0750 6.3450 0.0750 ;
        RECT 5.9250 -0.0750 6.0450 0.1950 ;
        RECT 5.6250 -0.0750 5.9250 0.0750 ;
        RECT 5.5050 -0.0750 5.6250 0.1950 ;
        RECT 5.2050 -0.0750 5.5050 0.0750 ;
        RECT 5.0850 -0.0750 5.2050 0.1950 ;
        RECT 4.7850 -0.0750 5.0850 0.0750 ;
        RECT 4.6650 -0.0750 4.7850 0.1950 ;
        RECT 4.3650 -0.0750 4.6650 0.0750 ;
        RECT 4.2450 -0.0750 4.3650 0.1950 ;
        RECT 3.9450 -0.0750 4.2450 0.0750 ;
        RECT 3.8250 -0.0750 3.9450 0.1950 ;
        RECT 3.5250 -0.0750 3.8250 0.0750 ;
        RECT 3.4050 -0.0750 3.5250 0.1950 ;
        RECT 3.1050 -0.0750 3.4050 0.0750 ;
        RECT 2.9850 -0.0750 3.1050 0.1950 ;
        RECT 2.6850 -0.0750 2.9850 0.0750 ;
        RECT 2.5650 -0.0750 2.6850 0.1950 ;
        RECT 2.2650 -0.0750 2.5650 0.0750 ;
        RECT 2.1450 -0.0750 2.2650 0.1950 ;
        RECT 1.8450 -0.0750 2.1450 0.0750 ;
        RECT 1.7250 -0.0750 1.8450 0.1950 ;
        RECT 1.4250 -0.0750 1.7250 0.0750 ;
        RECT 1.3050 -0.0750 1.4250 0.1950 ;
        RECT 1.0050 -0.0750 1.3050 0.0750 ;
        RECT 0.8850 -0.0750 1.0050 0.1950 ;
        RECT 0.5850 -0.0750 0.8850 0.0750 ;
        RECT 0.4650 -0.0750 0.5850 0.1950 ;
        RECT 0.1425 -0.0750 0.4650 0.0750 ;
        RECT 0.0675 -0.0750 0.1425 0.2625 ;
        RECT 0.0000 -0.0750 0.0675 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 6.6750 0.9750 6.9300 1.1250 ;
        RECT 6.5550 0.8250 6.6750 1.1250 ;
        RECT 6.2550 0.9750 6.5550 1.1250 ;
        RECT 6.1350 0.8250 6.2550 1.1250 ;
        RECT 5.8350 0.9750 6.1350 1.1250 ;
        RECT 5.7150 0.8250 5.8350 1.1250 ;
        RECT 5.4150 0.9750 5.7150 1.1250 ;
        RECT 5.2950 0.8250 5.4150 1.1250 ;
        RECT 4.9950 0.9750 5.2950 1.1250 ;
        RECT 4.8750 0.8250 4.9950 1.1250 ;
        RECT 4.5750 0.9750 4.8750 1.1250 ;
        RECT 4.4550 0.8250 4.5750 1.1250 ;
        RECT 4.1550 0.9750 4.4550 1.1250 ;
        RECT 4.0350 0.8250 4.1550 1.1250 ;
        RECT 3.7350 0.9750 4.0350 1.1250 ;
        RECT 3.6150 0.8250 3.7350 1.1250 ;
        RECT 0.0000 0.9750 3.6150 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 6.7950 0.1725 6.8550 0.2325 ;
        RECT 6.7950 0.6975 6.8550 0.7575 ;
        RECT 6.6900 0.4950 6.7500 0.5550 ;
        RECT 6.5850 0.3000 6.6450 0.3600 ;
        RECT 6.5850 0.8325 6.6450 0.8925 ;
        RECT 6.4800 0.4950 6.5400 0.5550 ;
        RECT 6.3750 0.1350 6.4350 0.1950 ;
        RECT 6.3750 0.6825 6.4350 0.7425 ;
        RECT 6.2700 0.4950 6.3300 0.5550 ;
        RECT 6.1650 0.3000 6.2250 0.3600 ;
        RECT 6.1650 0.8325 6.2250 0.8925 ;
        RECT 6.0600 0.4950 6.1200 0.5550 ;
        RECT 5.9550 0.1350 6.0150 0.1950 ;
        RECT 5.9550 0.6825 6.0150 0.7425 ;
        RECT 5.8500 0.4950 5.9100 0.5550 ;
        RECT 5.7450 0.3000 5.8050 0.3600 ;
        RECT 5.7450 0.8325 5.8050 0.8925 ;
        RECT 5.6400 0.4950 5.7000 0.5550 ;
        RECT 5.5350 0.1350 5.5950 0.1950 ;
        RECT 5.5350 0.6825 5.5950 0.7425 ;
        RECT 5.4300 0.4950 5.4900 0.5550 ;
        RECT 5.3250 0.3000 5.3850 0.3600 ;
        RECT 5.3250 0.8325 5.3850 0.8925 ;
        RECT 5.2200 0.4950 5.2800 0.5550 ;
        RECT 5.1150 0.1350 5.1750 0.1950 ;
        RECT 5.1150 0.6825 5.1750 0.7425 ;
        RECT 5.0100 0.4950 5.0700 0.5550 ;
        RECT 4.9050 0.3000 4.9650 0.3600 ;
        RECT 4.9050 0.8325 4.9650 0.8925 ;
        RECT 4.8000 0.4950 4.8600 0.5550 ;
        RECT 4.6950 0.1350 4.7550 0.1950 ;
        RECT 4.6950 0.6825 4.7550 0.7425 ;
        RECT 4.5900 0.4950 4.6500 0.5550 ;
        RECT 4.4850 0.3000 4.5450 0.3600 ;
        RECT 4.4850 0.8325 4.5450 0.8925 ;
        RECT 4.3800 0.4950 4.4400 0.5550 ;
        RECT 4.2750 0.1350 4.3350 0.1950 ;
        RECT 4.2750 0.6825 4.3350 0.7425 ;
        RECT 4.1700 0.4950 4.2300 0.5550 ;
        RECT 4.0650 0.3000 4.1250 0.3600 ;
        RECT 4.0650 0.8325 4.1250 0.8925 ;
        RECT 3.9600 0.4950 4.0200 0.5550 ;
        RECT 3.8550 0.1350 3.9150 0.1950 ;
        RECT 3.8550 0.6825 3.9150 0.7425 ;
        RECT 3.7500 0.4950 3.8100 0.5550 ;
        RECT 3.6450 0.3000 3.7050 0.3600 ;
        RECT 3.6450 0.8325 3.7050 0.8925 ;
        RECT 3.5400 0.4950 3.6000 0.5550 ;
        RECT 3.4350 0.1350 3.4950 0.1950 ;
        RECT 3.4350 0.7650 3.4950 0.8250 ;
        RECT 3.3300 0.4800 3.3900 0.5400 ;
        RECT 3.2250 0.3000 3.2850 0.3600 ;
        RECT 3.2250 0.6600 3.2850 0.7200 ;
        RECT 3.1200 0.4800 3.1800 0.5400 ;
        RECT 3.0150 0.1350 3.0750 0.1950 ;
        RECT 3.0150 0.8325 3.0750 0.8925 ;
        RECT 2.9100 0.4800 2.9700 0.5400 ;
        RECT 2.8050 0.3000 2.8650 0.3600 ;
        RECT 2.8050 0.6600 2.8650 0.7200 ;
        RECT 2.7000 0.4800 2.7600 0.5400 ;
        RECT 2.5950 0.1350 2.6550 0.1950 ;
        RECT 2.5950 0.8325 2.6550 0.8925 ;
        RECT 2.4900 0.4800 2.5500 0.5400 ;
        RECT 2.3850 0.3000 2.4450 0.3600 ;
        RECT 2.3850 0.6600 2.4450 0.7200 ;
        RECT 2.2800 0.4800 2.3400 0.5400 ;
        RECT 2.1750 0.1350 2.2350 0.1950 ;
        RECT 2.1750 0.8325 2.2350 0.8925 ;
        RECT 2.0700 0.4800 2.1300 0.5400 ;
        RECT 1.9650 0.3000 2.0250 0.3600 ;
        RECT 1.9650 0.6600 2.0250 0.7200 ;
        RECT 1.8600 0.4800 1.9200 0.5400 ;
        RECT 1.7550 0.1350 1.8150 0.1950 ;
        RECT 1.7550 0.8325 1.8150 0.8925 ;
        RECT 1.6500 0.4800 1.7100 0.5400 ;
        RECT 1.5450 0.3000 1.6050 0.3600 ;
        RECT 1.5450 0.6600 1.6050 0.7200 ;
        RECT 1.4400 0.4800 1.5000 0.5400 ;
        RECT 1.3350 0.1350 1.3950 0.1950 ;
        RECT 1.3350 0.8325 1.3950 0.8925 ;
        RECT 1.2300 0.4800 1.2900 0.5400 ;
        RECT 1.1250 0.3000 1.1850 0.3600 ;
        RECT 1.1250 0.6600 1.1850 0.7200 ;
        RECT 1.0200 0.4800 1.0800 0.5400 ;
        RECT 0.9150 0.1350 0.9750 0.1950 ;
        RECT 0.9150 0.8325 0.9750 0.8925 ;
        RECT 0.2850 0.3000 0.3450 0.3600 ;
        RECT 0.2850 0.6600 0.3450 0.7200 ;
        RECT 0.1800 0.4800 0.2400 0.5400 ;
        RECT 0.0750 0.1725 0.1350 0.2325 ;
        RECT 0.0750 0.8025 0.1350 0.8625 ;
        RECT 0.8100 0.4800 0.8700 0.5400 ;
        RECT 0.7050 0.3000 0.7650 0.3600 ;
        RECT 0.7050 0.6600 0.7650 0.7200 ;
        RECT 0.6000 0.4800 0.6600 0.5400 ;
        RECT 0.4950 0.1350 0.5550 0.1950 ;
        RECT 0.4950 0.8325 0.5550 0.8925 ;
        RECT 0.3900 0.4800 0.4500 0.5400 ;
        LAYER M1 ;
        RECT 6.7725 0.6750 6.8775 0.7800 ;
        RECT 3.5325 0.4650 6.7875 0.5850 ;
        RECT 3.5025 0.6750 6.7725 0.7500 ;
        RECT 0.2550 0.2700 6.6750 0.3900 ;
        RECT 3.4275 0.6750 3.5025 0.9000 ;
        RECT 0.1575 0.8250 3.4275 0.9000 ;
        RECT 0.2550 0.6300 3.3075 0.7500 ;
        RECT 0.0525 0.7800 0.1575 0.9000 ;
        LAYER M2 ;
        RECT 2.8125 0.2700 2.9400 0.3900 ;
        RECT 2.8125 0.6300 2.9400 0.7500 ;
        RECT 2.3100 0.2700 2.4375 0.3900 ;
        RECT 2.3100 0.6300 2.4375 0.7500 ;
    END
END NR2_1100


MACRO NR3_0001
    CLASS CORE ;
    FOREIGN NR3_0001 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.2000 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 0.7875 0.7125 1.3200 0.7875 ;
        RECT 0.6825 0.2475 0.7875 0.7875 ;
        VIA 0.7350 0.3300 VIA12_square ;
        VIA 0.7350 0.6975 VIA12_square ;
        END
    END ZN
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 3.2025 0.4125 3.3075 0.6000 ;
        RECT 2.7375 0.4125 3.2025 0.4875 ;
        VIA 3.2550 0.5175 VIA12_square ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 2.1525 0.4125 2.2575 0.6000 ;
        RECT 1.6875 0.4125 2.1525 0.4875 ;
        VIA 2.2050 0.5175 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1725 0.4650 1.3200 0.5700 ;
        RECT 0.0675 0.3675 0.1725 0.6825 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 4.1475 -0.0750 4.2000 0.0750 ;
        RECT 4.0425 -0.0750 4.1475 0.2625 ;
        RECT 3.7350 -0.0750 4.0425 0.0750 ;
        RECT 3.6150 -0.0750 3.7350 0.2175 ;
        RECT 3.3150 -0.0750 3.6150 0.0750 ;
        RECT 3.1950 -0.0750 3.3150 0.2175 ;
        RECT 2.8950 -0.0750 3.1950 0.0750 ;
        RECT 2.7750 -0.0750 2.8950 0.2175 ;
        RECT 2.6850 -0.0750 2.7750 0.0750 ;
        RECT 2.5650 -0.0750 2.6850 0.2175 ;
        RECT 2.2650 -0.0750 2.5650 0.0750 ;
        RECT 2.1450 -0.0750 2.2650 0.2175 ;
        RECT 1.8450 -0.0750 2.1450 0.0750 ;
        RECT 1.7250 -0.0750 1.8450 0.2175 ;
        RECT 1.4250 -0.0750 1.7250 0.0750 ;
        RECT 1.3050 -0.0750 1.4250 0.2175 ;
        RECT 1.0050 -0.0750 1.3050 0.0750 ;
        RECT 0.8850 -0.0750 1.0050 0.2175 ;
        RECT 0.5850 -0.0750 0.8850 0.0750 ;
        RECT 0.4650 -0.0750 0.5850 0.2175 ;
        RECT 0.1425 -0.0750 0.4650 0.0750 ;
        RECT 0.0675 -0.0750 0.1425 0.2475 ;
        RECT 0.0000 -0.0750 0.0675 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 3.9450 0.9750 4.2000 1.1250 ;
        RECT 3.8250 0.8175 3.9450 1.1250 ;
        RECT 3.5250 0.9750 3.8250 1.1250 ;
        RECT 3.4050 0.8175 3.5250 1.1250 ;
        RECT 3.1050 0.9750 3.4050 1.1250 ;
        RECT 2.9850 0.8175 3.1050 1.1250 ;
        RECT 0.0000 0.9750 2.9850 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 4.0650 0.1575 4.1250 0.2175 ;
        RECT 4.0650 0.7350 4.1250 0.7950 ;
        RECT 3.9600 0.4875 4.0200 0.5475 ;
        RECT 3.8550 0.1575 3.9150 0.2175 ;
        RECT 3.8550 0.8400 3.9150 0.9000 ;
        RECT 3.7500 0.4875 3.8100 0.5475 ;
        RECT 3.6450 0.1425 3.7050 0.2025 ;
        RECT 3.6450 0.6750 3.7050 0.7350 ;
        RECT 3.5400 0.4875 3.6000 0.5475 ;
        RECT 3.4350 0.1575 3.4950 0.2175 ;
        RECT 3.4350 0.8400 3.4950 0.9000 ;
        RECT 3.3300 0.4875 3.3900 0.5475 ;
        RECT 3.2250 0.1425 3.2850 0.2025 ;
        RECT 3.2250 0.6750 3.2850 0.7350 ;
        RECT 3.1200 0.4875 3.1800 0.5475 ;
        RECT 3.0150 0.1575 3.0750 0.2175 ;
        RECT 3.0150 0.8400 3.0750 0.9000 ;
        RECT 2.9100 0.4875 2.9700 0.5475 ;
        RECT 2.8050 0.1575 2.8650 0.2175 ;
        RECT 2.8050 0.6750 2.8650 0.7350 ;
        RECT 2.5950 0.1575 2.6550 0.2175 ;
        RECT 2.5950 0.8325 2.6550 0.8925 ;
        RECT 2.4900 0.4875 2.5500 0.5475 ;
        RECT 2.3850 0.1575 2.4450 0.2175 ;
        RECT 2.3850 0.6750 2.4450 0.7350 ;
        RECT 2.2800 0.4875 2.3400 0.5475 ;
        RECT 2.1750 0.1425 2.2350 0.2025 ;
        RECT 2.1750 0.8325 2.2350 0.8925 ;
        RECT 2.0700 0.4875 2.1300 0.5475 ;
        RECT 1.9650 0.1575 2.0250 0.2175 ;
        RECT 1.9650 0.6750 2.0250 0.7350 ;
        RECT 1.8600 0.4875 1.9200 0.5475 ;
        RECT 1.7550 0.1425 1.8150 0.2025 ;
        RECT 1.7550 0.8325 1.8150 0.8925 ;
        RECT 1.6500 0.4875 1.7100 0.5475 ;
        RECT 1.5450 0.1575 1.6050 0.2175 ;
        RECT 1.5450 0.6750 1.6050 0.7350 ;
        RECT 1.4400 0.4875 1.5000 0.5475 ;
        RECT 1.3350 0.1425 1.3950 0.2025 ;
        RECT 1.3350 0.8325 1.3950 0.8925 ;
        RECT 1.2300 0.4875 1.2900 0.5475 ;
        RECT 1.1250 0.1575 1.1850 0.2175 ;
        RECT 1.1250 0.6675 1.1850 0.7275 ;
        RECT 1.0200 0.4875 1.0800 0.5475 ;
        RECT 0.9150 0.1425 0.9750 0.2025 ;
        RECT 0.9150 0.8325 0.9750 0.8925 ;
        RECT 0.8100 0.4875 0.8700 0.5475 ;
        RECT 0.7050 0.1575 0.7650 0.2175 ;
        RECT 0.7050 0.6675 0.7650 0.7275 ;
        RECT 0.6000 0.4875 0.6600 0.5475 ;
        RECT 0.4950 0.1425 0.5550 0.2025 ;
        RECT 0.4950 0.8325 0.5550 0.8925 ;
        RECT 0.3900 0.4875 0.4500 0.5475 ;
        RECT 0.2850 0.1575 0.3450 0.2175 ;
        RECT 0.2850 0.6675 0.3450 0.7275 ;
        RECT 0.1800 0.4875 0.2400 0.5475 ;
        RECT 0.0750 0.1575 0.1350 0.2175 ;
        RECT 0.0750 0.8025 0.1350 0.8625 ;
        LAYER M1 ;
        RECT 4.0575 0.6675 4.1325 0.8250 ;
        RECT 2.8800 0.4650 4.0650 0.5700 ;
        RECT 1.5000 0.6675 4.0575 0.7425 ;
        RECT 3.8250 0.1500 3.9450 0.3675 ;
        RECT 3.5250 0.2925 3.8250 0.3675 ;
        RECT 3.4050 0.1500 3.5250 0.3675 ;
        RECT 3.1050 0.2925 3.4050 0.3675 ;
        RECT 2.9850 0.1500 3.1050 0.3675 ;
        RECT 2.4750 0.2925 2.9850 0.3675 ;
        RECT 0.1575 0.8250 2.7000 0.9000 ;
        RECT 1.4175 0.4650 2.6100 0.5700 ;
        RECT 2.3550 0.1500 2.4750 0.3675 ;
        RECT 2.0550 0.2925 2.3550 0.3675 ;
        RECT 1.9350 0.1500 2.0550 0.3675 ;
        RECT 1.6350 0.2925 1.9350 0.3675 ;
        RECT 1.5150 0.1500 1.6350 0.3675 ;
        RECT 1.2150 0.2925 1.5150 0.3675 ;
        RECT 1.0950 0.1500 1.2150 0.3675 ;
        RECT 0.2625 0.6450 1.2150 0.7500 ;
        RECT 0.7950 0.2925 1.0950 0.3675 ;
        RECT 0.6750 0.1500 0.7950 0.3675 ;
        RECT 0.3750 0.2925 0.6750 0.3675 ;
        RECT 0.2550 0.1500 0.3750 0.3675 ;
        RECT 0.0525 0.7725 0.1575 0.9000 ;
    END
END NR3_0001


MACRO NR3_0010
    CLASS CORE ;
    FOREIGN NR3_0010 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.7200 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 1.3125 0.3000 1.4700 0.4200 ;
        RECT 1.3125 0.6375 1.4700 0.7575 ;
        RECT 0.9975 0.3000 1.3125 0.7575 ;
        RECT 0.8400 0.3000 0.9975 0.4200 ;
        RECT 0.8400 0.6375 0.9975 0.7575 ;
        VIA 1.3125 0.3600 VIA12_slot ;
        VIA 1.3125 0.6975 VIA12_slot ;
        VIA 0.9975 0.3600 VIA12_slot ;
        VIA 0.9975 0.6975 VIA12_slot ;
        END
    END ZN
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 6.5325 0.3675 6.6375 0.6375 ;
        RECT 6.4725 0.4950 6.5325 0.6375 ;
        RECT 4.1400 0.4950 6.4725 0.5700 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 2.2575 0.4500 2.3625 0.6375 ;
        RECT 1.8975 0.5625 2.2575 0.6375 ;
        VIA 2.3100 0.5475 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1425 0.4950 1.7400 0.5700 ;
        RECT 0.0675 0.3675 0.1425 0.6825 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 6.6525 -0.0750 6.7200 0.0750 ;
        RECT 6.5775 -0.0750 6.6525 0.2625 ;
        RECT 6.2475 -0.0750 6.5775 0.0750 ;
        RECT 6.1425 -0.0750 6.2475 0.2250 ;
        RECT 5.8275 -0.0750 6.1425 0.0750 ;
        RECT 5.7225 -0.0750 5.8275 0.2250 ;
        RECT 5.4075 -0.0750 5.7225 0.0750 ;
        RECT 5.3025 -0.0750 5.4075 0.2250 ;
        RECT 4.9875 -0.0750 5.3025 0.0750 ;
        RECT 4.8825 -0.0750 4.9875 0.2250 ;
        RECT 4.5675 -0.0750 4.8825 0.0750 ;
        RECT 4.4625 -0.0750 4.5675 0.2250 ;
        RECT 4.1550 -0.0750 4.4625 0.0750 ;
        RECT 4.0350 -0.0750 4.1550 0.2250 ;
        RECT 3.9450 -0.0750 4.0350 0.0750 ;
        RECT 3.8250 -0.0750 3.9450 0.2250 ;
        RECT 3.5250 -0.0750 3.8250 0.0750 ;
        RECT 3.4050 -0.0750 3.5250 0.2250 ;
        RECT 3.0975 -0.0750 3.4050 0.0750 ;
        RECT 2.9925 -0.0750 3.0975 0.2250 ;
        RECT 2.6775 -0.0750 2.9925 0.0750 ;
        RECT 2.5725 -0.0750 2.6775 0.2250 ;
        RECT 2.2650 -0.0750 2.5725 0.0750 ;
        RECT 2.1450 -0.0750 2.2650 0.1950 ;
        RECT 1.8450 -0.0750 2.1450 0.0750 ;
        RECT 1.7250 -0.0750 1.8450 0.1950 ;
        RECT 1.4175 -0.0750 1.7250 0.0750 ;
        RECT 1.3125 -0.0750 1.4175 0.2250 ;
        RECT 0.9975 -0.0750 1.3125 0.0750 ;
        RECT 0.8925 -0.0750 0.9975 0.2250 ;
        RECT 0.5775 -0.0750 0.8925 0.0750 ;
        RECT 0.4725 -0.0750 0.5775 0.2250 ;
        RECT 0.1425 -0.0750 0.4725 0.0750 ;
        RECT 0.0675 -0.0750 0.1425 0.2475 ;
        RECT 0.0000 -0.0750 0.0675 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 6.4650 0.9750 6.7200 1.1250 ;
        RECT 6.3450 0.8625 6.4650 1.1250 ;
        RECT 6.0450 0.9750 6.3450 1.1250 ;
        RECT 5.9250 0.8400 6.0450 1.1250 ;
        RECT 5.6250 0.9750 5.9250 1.1250 ;
        RECT 5.5050 0.8400 5.6250 1.1250 ;
        RECT 5.2050 0.9750 5.5050 1.1250 ;
        RECT 5.0850 0.8400 5.2050 1.1250 ;
        RECT 4.7850 0.9750 5.0850 1.1250 ;
        RECT 4.6650 0.8400 4.7850 1.1250 ;
        RECT 4.3650 0.9750 4.6650 1.1250 ;
        RECT 4.2450 0.8400 4.3650 1.1250 ;
        RECT 0.0000 0.9750 4.2450 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 6.5850 0.1575 6.6450 0.2175 ;
        RECT 6.5850 0.7800 6.6450 0.8400 ;
        RECT 6.4800 0.4950 6.5400 0.5550 ;
        RECT 6.3750 0.1725 6.4350 0.2325 ;
        RECT 6.3750 0.8625 6.4350 0.9225 ;
        RECT 6.2700 0.4950 6.3300 0.5550 ;
        RECT 6.1650 0.1350 6.2250 0.1950 ;
        RECT 6.1650 0.6900 6.2250 0.7500 ;
        RECT 6.0600 0.4950 6.1200 0.5550 ;
        RECT 5.9550 0.1725 6.0150 0.2325 ;
        RECT 5.9550 0.8550 6.0150 0.9150 ;
        RECT 5.8500 0.4950 5.9100 0.5550 ;
        RECT 5.7450 0.1350 5.8050 0.1950 ;
        RECT 5.7450 0.6900 5.8050 0.7500 ;
        RECT 5.6400 0.4950 5.7000 0.5550 ;
        RECT 5.5350 0.1725 5.5950 0.2325 ;
        RECT 5.5350 0.8550 5.5950 0.9150 ;
        RECT 5.4300 0.4950 5.4900 0.5550 ;
        RECT 5.3250 0.1350 5.3850 0.1950 ;
        RECT 5.3250 0.6900 5.3850 0.7500 ;
        RECT 5.2200 0.4950 5.2800 0.5550 ;
        RECT 5.1150 0.1725 5.1750 0.2325 ;
        RECT 5.1150 0.8550 5.1750 0.9150 ;
        RECT 5.0100 0.4950 5.0700 0.5550 ;
        RECT 4.9050 0.1350 4.9650 0.1950 ;
        RECT 4.9050 0.6900 4.9650 0.7500 ;
        RECT 4.8000 0.4950 4.8600 0.5550 ;
        RECT 4.6950 0.3225 4.7550 0.3825 ;
        RECT 4.6950 0.8550 4.7550 0.9150 ;
        RECT 4.5900 0.4950 4.6500 0.5550 ;
        RECT 4.4850 0.1350 4.5450 0.1950 ;
        RECT 4.4850 0.6900 4.5450 0.7500 ;
        RECT 4.3800 0.4950 4.4400 0.5550 ;
        RECT 4.2750 0.3225 4.3350 0.3825 ;
        RECT 4.2750 0.8550 4.3350 0.9150 ;
        RECT 4.1700 0.4950 4.2300 0.5550 ;
        RECT 4.0650 0.1575 4.1250 0.2175 ;
        RECT 4.0650 0.6900 4.1250 0.7500 ;
        RECT 3.8550 0.1575 3.9150 0.2175 ;
        RECT 3.8550 0.8325 3.9150 0.8925 ;
        RECT 3.7500 0.4950 3.8100 0.5550 ;
        RECT 3.6450 0.1725 3.7050 0.2325 ;
        RECT 3.6450 0.6900 3.7050 0.7500 ;
        RECT 3.5400 0.4950 3.6000 0.5550 ;
        RECT 3.4350 0.1575 3.4950 0.2175 ;
        RECT 3.4350 0.8325 3.4950 0.8925 ;
        RECT 3.3300 0.4950 3.3900 0.5550 ;
        RECT 3.2250 0.1725 3.2850 0.2325 ;
        RECT 3.2250 0.6900 3.2850 0.7500 ;
        RECT 3.1200 0.4950 3.1800 0.5550 ;
        RECT 3.0150 0.1350 3.0750 0.1950 ;
        RECT 3.0150 0.8325 3.0750 0.8925 ;
        RECT 2.9100 0.4950 2.9700 0.5550 ;
        RECT 2.8050 0.3225 2.8650 0.3825 ;
        RECT 2.8050 0.6900 2.8650 0.7500 ;
        RECT 2.7000 0.4950 2.7600 0.5550 ;
        RECT 2.5950 0.1350 2.6550 0.1950 ;
        RECT 2.5950 0.8325 2.6550 0.8925 ;
        RECT 2.4900 0.4950 2.5500 0.5550 ;
        RECT 2.3850 0.3225 2.4450 0.3825 ;
        RECT 2.3850 0.6900 2.4450 0.7500 ;
        RECT 2.2800 0.4950 2.3400 0.5550 ;
        RECT 2.1750 0.1350 2.2350 0.1950 ;
        RECT 2.1750 0.8325 2.2350 0.8925 ;
        RECT 2.0700 0.4950 2.1300 0.5550 ;
        RECT 1.9650 0.3225 2.0250 0.3825 ;
        RECT 1.9650 0.6900 2.0250 0.7500 ;
        RECT 1.8600 0.4950 1.9200 0.5550 ;
        RECT 1.7550 0.1350 1.8150 0.1950 ;
        RECT 1.7550 0.8325 1.8150 0.8925 ;
        RECT 1.6500 0.4950 1.7100 0.5550 ;
        RECT 1.5450 0.3225 1.6050 0.3825 ;
        RECT 1.5450 0.6900 1.6050 0.7500 ;
        RECT 1.4400 0.4950 1.5000 0.5550 ;
        RECT 1.3350 0.1350 1.3950 0.1950 ;
        RECT 1.3350 0.8325 1.3950 0.8925 ;
        RECT 1.2300 0.4950 1.2900 0.5550 ;
        RECT 1.1250 0.3225 1.1850 0.3825 ;
        RECT 1.1250 0.6900 1.1850 0.7500 ;
        RECT 1.0200 0.4950 1.0800 0.5550 ;
        RECT 0.9150 0.1350 0.9750 0.1950 ;
        RECT 0.9150 0.8325 0.9750 0.8925 ;
        RECT 0.8100 0.4950 0.8700 0.5550 ;
        RECT 0.7050 0.3225 0.7650 0.3825 ;
        RECT 0.7050 0.6900 0.7650 0.7500 ;
        RECT 0.6000 0.4950 0.6600 0.5550 ;
        RECT 0.4950 0.1350 0.5550 0.1950 ;
        RECT 0.4950 0.8325 0.5550 0.8925 ;
        RECT 0.3900 0.4950 0.4500 0.5550 ;
        RECT 0.2850 0.3225 0.3450 0.3825 ;
        RECT 0.2850 0.6900 0.3450 0.7500 ;
        RECT 0.1800 0.4950 0.2400 0.5550 ;
        RECT 0.0750 0.1575 0.1350 0.2175 ;
        RECT 0.0750 0.8175 0.1350 0.8775 ;
        LAYER M1 ;
        RECT 6.5775 0.7125 6.6525 0.8700 ;
        RECT 6.3975 0.7125 6.5775 0.7875 ;
        RECT 6.3525 0.1500 6.4575 0.4200 ;
        RECT 6.3225 0.6750 6.3975 0.7875 ;
        RECT 6.0375 0.3000 6.3525 0.4200 ;
        RECT 1.9350 0.6750 6.3225 0.7500 ;
        RECT 5.9325 0.1500 6.0375 0.4200 ;
        RECT 5.6175 0.3000 5.9325 0.4200 ;
        RECT 5.5125 0.1500 5.6175 0.4200 ;
        RECT 5.1975 0.3000 5.5125 0.4200 ;
        RECT 5.0925 0.1500 5.1975 0.4200 ;
        RECT 3.7275 0.3000 5.0925 0.4200 ;
        RECT 0.1575 0.8250 3.9600 0.9000 ;
        RECT 1.9650 0.4950 3.8625 0.6000 ;
        RECT 3.6225 0.1500 3.7275 0.4200 ;
        RECT 3.3075 0.3000 3.6225 0.4200 ;
        RECT 3.2025 0.1500 3.3075 0.4200 ;
        RECT 2.1675 0.3000 3.2025 0.4200 ;
        RECT 2.0475 0.2700 2.1675 0.4200 ;
        RECT 1.7850 0.2700 2.0475 0.3900 ;
        RECT 1.8600 0.4650 1.9650 0.6000 ;
        RECT 1.6650 0.2700 1.7850 0.4200 ;
        RECT 0.2550 0.3000 1.6650 0.4200 ;
        RECT 0.2550 0.6450 1.6500 0.7500 ;
        RECT 0.0525 0.7950 0.1575 0.9000 ;
        LAYER M2 ;
        RECT 1.3425 0.3000 1.4700 0.4200 ;
        RECT 1.3425 0.6375 1.4700 0.7575 ;
        RECT 0.8400 0.3000 0.9675 0.4200 ;
        RECT 0.8400 0.6375 0.9675 0.7575 ;
    END
END NR3_0010


MACRO NR3_0011
    CLASS CORE ;
    FOREIGN NR3_0011 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.4700 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 0.9675 0.8625 1.2825 0.9375 ;
        RECT 0.8925 0.2625 0.9675 0.9375 ;
        RECT 0.5775 0.2625 0.8925 0.3375 ;
        RECT 0.5025 0.2625 0.5775 0.3675 ;
        VIA 0.9300 0.8325 VIA12_square ;
        VIA 0.8100 0.3000 VIA12_square ;
        END
    END ZN
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.2300 0.4200 1.3350 0.7200 ;
        RECT 0.1425 0.6450 1.2300 0.7200 ;
        RECT 0.1425 0.4200 0.2325 0.5550 ;
        RECT 0.0675 0.3675 0.1425 0.7200 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.0425 0.1125 1.1175 0.6450 ;
        RECT 0.4275 0.1125 1.0425 0.1875 ;
        RECT 0.3525 0.1125 0.4275 0.5400 ;
        VIA 1.0800 0.4950 VIA12_square ;
        VIA 0.3900 0.4575 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.6825 0.4125 0.7875 0.7875 ;
        RECT 0.2175 0.7125 0.6825 0.7875 ;
        VIA 0.7350 0.4950 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.4250 -0.0750 1.4700 0.0750 ;
        RECT 1.3050 -0.0750 1.4250 0.2475 ;
        RECT 1.0050 -0.0750 1.3050 0.0750 ;
        RECT 0.8850 -0.0750 1.0050 0.1875 ;
        RECT 0.5850 -0.0750 0.8850 0.0750 ;
        RECT 0.4650 -0.0750 0.5850 0.1875 ;
        RECT 0.1650 -0.0750 0.4650 0.0750 ;
        RECT 0.0450 -0.0750 0.1650 0.2475 ;
        RECT 0.0000 -0.0750 0.0450 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.4175 0.9750 1.4700 1.1250 ;
        RECT 1.3125 0.8100 1.4175 1.1250 ;
        RECT 0.1575 0.9750 1.3125 1.1250 ;
        RECT 0.0525 0.8100 0.1575 1.1250 ;
        RECT 0.0000 0.9750 0.0525 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.3350 0.1575 1.3950 0.2175 ;
        RECT 1.3350 0.8325 1.3950 0.8925 ;
        RECT 1.2300 0.4650 1.2900 0.5250 ;
        RECT 1.1250 0.1800 1.1850 0.2400 ;
        RECT 1.0200 0.4650 1.0800 0.5250 ;
        RECT 0.9150 0.1275 0.9750 0.1875 ;
        RECT 0.8100 0.4650 0.8700 0.5250 ;
        RECT 0.7050 0.1800 0.7650 0.2400 ;
        RECT 0.7050 0.8025 0.7650 0.8625 ;
        RECT 0.6000 0.4650 0.6600 0.5250 ;
        RECT 0.4950 0.1275 0.5550 0.1875 ;
        RECT 0.3900 0.4650 0.4500 0.5250 ;
        RECT 0.2850 0.1800 0.3450 0.2400 ;
        RECT 0.1725 0.4650 0.2325 0.5250 ;
        RECT 0.0750 0.1575 0.1350 0.2175 ;
        RECT 0.0750 0.8325 0.1350 0.8925 ;
        LAYER M1 ;
        RECT 1.1025 0.1575 1.2075 0.3375 ;
        RECT 0.9450 0.4200 1.1550 0.5700 ;
        RECT 0.7875 0.2625 1.1025 0.3375 ;
        RECT 0.6000 0.7950 1.0650 0.8700 ;
        RECT 0.6825 0.1575 0.7875 0.3375 ;
        RECT 0.3675 0.2625 0.6825 0.3375 ;
        RECT 0.3075 0.4200 0.5250 0.5700 ;
        RECT 0.2625 0.1575 0.3675 0.3375 ;
        RECT 0.6000 0.4350 0.8700 0.5550 ;
    END
END NR3_0011


MACRO NR3_0100
    CLASS CORE ;
    FOREIGN NR3_0100 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.5000 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 1.9425 0.2775 2.1000 0.3975 ;
        RECT 1.9425 0.6375 2.1000 0.7575 ;
        RECT 1.6275 0.2775 1.9425 0.7575 ;
        RECT 1.4700 0.2775 1.6275 0.3975 ;
        RECT 1.4700 0.6375 1.6275 0.7575 ;
        VIA 1.9425 0.3375 VIA12_slot ;
        VIA 1.9425 0.6975 VIA12_slot ;
        VIA 1.6275 0.3375 VIA12_slot ;
        VIA 1.6275 0.6975 VIA12_slot ;
        END
    END ZN
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 7.6125 0.4125 7.7175 0.6000 ;
        RECT 7.1475 0.4125 7.6125 0.4875 ;
        VIA 7.6650 0.5175 VIA12_square ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 4.2525 0.4125 4.3575 0.6000 ;
        RECT 3.7875 0.4125 4.2525 0.4875 ;
        VIA 4.3050 0.5175 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1725 0.4650 3.4200 0.5700 ;
        RECT 0.0675 0.3675 0.1725 0.6825 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 10.4475 -0.0750 10.5000 0.0750 ;
        RECT 10.3425 -0.0750 10.4475 0.2625 ;
        RECT 10.0350 -0.0750 10.3425 0.0750 ;
        RECT 9.9150 -0.0750 10.0350 0.2175 ;
        RECT 9.6150 -0.0750 9.9150 0.0750 ;
        RECT 9.4950 -0.0750 9.6150 0.2175 ;
        RECT 9.1950 -0.0750 9.4950 0.0750 ;
        RECT 9.0750 -0.0750 9.1950 0.2175 ;
        RECT 8.7750 -0.0750 9.0750 0.0750 ;
        RECT 8.6550 -0.0750 8.7750 0.2175 ;
        RECT 8.3550 -0.0750 8.6550 0.0750 ;
        RECT 8.2350 -0.0750 8.3550 0.2175 ;
        RECT 7.9350 -0.0750 8.2350 0.0750 ;
        RECT 7.8150 -0.0750 7.9350 0.2175 ;
        RECT 7.5150 -0.0750 7.8150 0.0750 ;
        RECT 7.3950 -0.0750 7.5150 0.2175 ;
        RECT 7.0950 -0.0750 7.3950 0.0750 ;
        RECT 6.9750 -0.0750 7.0950 0.2175 ;
        RECT 6.8850 -0.0750 6.9750 0.0750 ;
        RECT 6.7650 -0.0750 6.8850 0.2175 ;
        RECT 6.4650 -0.0750 6.7650 0.0750 ;
        RECT 6.3450 -0.0750 6.4650 0.2175 ;
        RECT 6.0450 -0.0750 6.3450 0.0750 ;
        RECT 5.9250 -0.0750 6.0450 0.2175 ;
        RECT 5.6250 -0.0750 5.9250 0.0750 ;
        RECT 5.5050 -0.0750 5.6250 0.2175 ;
        RECT 5.2050 -0.0750 5.5050 0.0750 ;
        RECT 5.0850 -0.0750 5.2050 0.2175 ;
        RECT 4.7850 -0.0750 5.0850 0.0750 ;
        RECT 4.6650 -0.0750 4.7850 0.2175 ;
        RECT 4.3650 -0.0750 4.6650 0.0750 ;
        RECT 4.2450 -0.0750 4.3650 0.2175 ;
        RECT 3.9450 -0.0750 4.2450 0.0750 ;
        RECT 3.8250 -0.0750 3.9450 0.2175 ;
        RECT 3.5250 -0.0750 3.8250 0.0750 ;
        RECT 3.4050 -0.0750 3.5250 0.2175 ;
        RECT 3.1050 -0.0750 3.4050 0.0750 ;
        RECT 2.9850 -0.0750 3.1050 0.2175 ;
        RECT 2.6850 -0.0750 2.9850 0.0750 ;
        RECT 2.5650 -0.0750 2.6850 0.2175 ;
        RECT 2.2650 -0.0750 2.5650 0.0750 ;
        RECT 2.1450 -0.0750 2.2650 0.2175 ;
        RECT 1.8450 -0.0750 2.1450 0.0750 ;
        RECT 1.7250 -0.0750 1.8450 0.2175 ;
        RECT 1.4250 -0.0750 1.7250 0.0750 ;
        RECT 1.3050 -0.0750 1.4250 0.2175 ;
        RECT 1.0050 -0.0750 1.3050 0.0750 ;
        RECT 0.8850 -0.0750 1.0050 0.2175 ;
        RECT 0.5850 -0.0750 0.8850 0.0750 ;
        RECT 0.4650 -0.0750 0.5850 0.2175 ;
        RECT 0.1425 -0.0750 0.4650 0.0750 ;
        RECT 0.0675 -0.0750 0.1425 0.2475 ;
        RECT 0.0000 -0.0750 0.0675 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 10.2450 0.9750 10.5000 1.1250 ;
        RECT 10.1250 0.8175 10.2450 1.1250 ;
        RECT 9.8250 0.9750 10.1250 1.1250 ;
        RECT 9.7050 0.8175 9.8250 1.1250 ;
        RECT 9.4050 0.9750 9.7050 1.1250 ;
        RECT 9.2850 0.8175 9.4050 1.1250 ;
        RECT 8.9850 0.9750 9.2850 1.1250 ;
        RECT 8.8650 0.8175 8.9850 1.1250 ;
        RECT 8.5650 0.9750 8.8650 1.1250 ;
        RECT 8.4450 0.8175 8.5650 1.1250 ;
        RECT 8.1450 0.9750 8.4450 1.1250 ;
        RECT 8.0250 0.8175 8.1450 1.1250 ;
        RECT 7.7250 0.9750 8.0250 1.1250 ;
        RECT 7.6050 0.8175 7.7250 1.1250 ;
        RECT 7.3050 0.9750 7.6050 1.1250 ;
        RECT 7.1850 0.8175 7.3050 1.1250 ;
        RECT 0.0000 0.9750 7.1850 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 10.3650 0.1575 10.4250 0.2175 ;
        RECT 10.3650 0.7350 10.4250 0.7950 ;
        RECT 10.2600 0.4875 10.3200 0.5475 ;
        RECT 10.1550 0.1725 10.2150 0.2325 ;
        RECT 10.1550 0.8400 10.2150 0.9000 ;
        RECT 10.0500 0.4875 10.1100 0.5475 ;
        RECT 9.9450 0.1425 10.0050 0.2025 ;
        RECT 9.9450 0.6750 10.0050 0.7350 ;
        RECT 9.8400 0.4875 9.9000 0.5475 ;
        RECT 9.7350 0.1725 9.7950 0.2325 ;
        RECT 9.7350 0.8400 9.7950 0.9000 ;
        RECT 9.6300 0.4875 9.6900 0.5475 ;
        RECT 9.5250 0.1425 9.5850 0.2025 ;
        RECT 9.5250 0.6750 9.5850 0.7350 ;
        RECT 9.4200 0.4875 9.4800 0.5475 ;
        RECT 9.3150 0.1725 9.3750 0.2325 ;
        RECT 9.3150 0.8400 9.3750 0.9000 ;
        RECT 9.2100 0.4875 9.2700 0.5475 ;
        RECT 9.1050 0.1425 9.1650 0.2025 ;
        RECT 9.1050 0.6750 9.1650 0.7350 ;
        RECT 9.0000 0.4875 9.0600 0.5475 ;
        RECT 8.8950 0.1725 8.9550 0.2325 ;
        RECT 8.8950 0.8400 8.9550 0.9000 ;
        RECT 8.7900 0.4875 8.8500 0.5475 ;
        RECT 8.6850 0.1425 8.7450 0.2025 ;
        RECT 8.6850 0.6750 8.7450 0.7350 ;
        RECT 8.5800 0.4875 8.6400 0.5475 ;
        RECT 8.4750 0.1725 8.5350 0.2325 ;
        RECT 8.4750 0.8400 8.5350 0.9000 ;
        RECT 8.3700 0.4875 8.4300 0.5475 ;
        RECT 8.2650 0.1425 8.3250 0.2025 ;
        RECT 8.2650 0.6750 8.3250 0.7350 ;
        RECT 8.1600 0.4875 8.2200 0.5475 ;
        RECT 8.0550 0.1575 8.1150 0.2175 ;
        RECT 8.0550 0.8400 8.1150 0.9000 ;
        RECT 7.9500 0.4875 8.0100 0.5475 ;
        RECT 7.8450 0.1425 7.9050 0.2025 ;
        RECT 7.8450 0.6750 7.9050 0.7350 ;
        RECT 7.7400 0.4875 7.8000 0.5475 ;
        RECT 7.6350 0.1575 7.6950 0.2175 ;
        RECT 7.6350 0.8400 7.6950 0.9000 ;
        RECT 7.5300 0.4875 7.5900 0.5475 ;
        RECT 7.4250 0.1425 7.4850 0.2025 ;
        RECT 7.4250 0.6750 7.4850 0.7350 ;
        RECT 7.3200 0.4875 7.3800 0.5475 ;
        RECT 7.2150 0.1575 7.2750 0.2175 ;
        RECT 7.2150 0.8400 7.2750 0.9000 ;
        RECT 7.1100 0.4875 7.1700 0.5475 ;
        RECT 7.0050 0.1575 7.0650 0.2175 ;
        RECT 7.0050 0.6750 7.0650 0.7350 ;
        RECT 6.7950 0.1575 6.8550 0.2175 ;
        RECT 6.7950 0.8325 6.8550 0.8925 ;
        RECT 6.6900 0.4875 6.7500 0.5475 ;
        RECT 6.5850 0.1575 6.6450 0.2175 ;
        RECT 6.5850 0.6750 6.6450 0.7350 ;
        RECT 6.4800 0.4875 6.5400 0.5475 ;
        RECT 6.3750 0.1425 6.4350 0.2025 ;
        RECT 6.3750 0.8325 6.4350 0.8925 ;
        RECT 6.2700 0.4875 6.3300 0.5475 ;
        RECT 6.1650 0.1575 6.2250 0.2175 ;
        RECT 6.1650 0.6750 6.2250 0.7350 ;
        RECT 6.0600 0.4875 6.1200 0.5475 ;
        RECT 5.9550 0.1425 6.0150 0.2025 ;
        RECT 5.9550 0.8325 6.0150 0.8925 ;
        RECT 5.8500 0.4875 5.9100 0.5475 ;
        RECT 5.7450 0.1575 5.8050 0.2175 ;
        RECT 5.7450 0.6750 5.8050 0.7350 ;
        RECT 5.6400 0.4875 5.7000 0.5475 ;
        RECT 5.5350 0.1425 5.5950 0.2025 ;
        RECT 5.5350 0.8325 5.5950 0.8925 ;
        RECT 5.4300 0.4875 5.4900 0.5475 ;
        RECT 5.3250 0.1575 5.3850 0.2175 ;
        RECT 5.3250 0.6750 5.3850 0.7350 ;
        RECT 5.2200 0.4875 5.2800 0.5475 ;
        RECT 5.1150 0.1425 5.1750 0.2025 ;
        RECT 5.1150 0.8325 5.1750 0.8925 ;
        RECT 5.0100 0.4875 5.0700 0.5475 ;
        RECT 4.9050 0.1575 4.9650 0.2175 ;
        RECT 4.9050 0.6750 4.9650 0.7350 ;
        RECT 4.8000 0.4875 4.8600 0.5475 ;
        RECT 4.6950 0.1425 4.7550 0.2025 ;
        RECT 4.6950 0.8325 4.7550 0.8925 ;
        RECT 4.5900 0.4875 4.6500 0.5475 ;
        RECT 4.4850 0.1575 4.5450 0.2175 ;
        RECT 4.4850 0.6750 4.5450 0.7350 ;
        RECT 4.3800 0.4875 4.4400 0.5475 ;
        RECT 4.2750 0.1425 4.3350 0.2025 ;
        RECT 4.2750 0.8325 4.3350 0.8925 ;
        RECT 4.1700 0.4875 4.2300 0.5475 ;
        RECT 4.0650 0.1575 4.1250 0.2175 ;
        RECT 4.0650 0.6750 4.1250 0.7350 ;
        RECT 3.9600 0.4875 4.0200 0.5475 ;
        RECT 3.8550 0.1425 3.9150 0.2025 ;
        RECT 3.8550 0.8325 3.9150 0.8925 ;
        RECT 3.7500 0.4875 3.8100 0.5475 ;
        RECT 3.6450 0.1575 3.7050 0.2175 ;
        RECT 3.6450 0.6750 3.7050 0.7350 ;
        RECT 3.5400 0.4875 3.6000 0.5475 ;
        RECT 3.4350 0.1425 3.4950 0.2025 ;
        RECT 3.4350 0.8325 3.4950 0.8925 ;
        RECT 3.3300 0.4875 3.3900 0.5475 ;
        RECT 3.2250 0.1575 3.2850 0.2175 ;
        RECT 3.2250 0.6675 3.2850 0.7275 ;
        RECT 3.1200 0.4875 3.1800 0.5475 ;
        RECT 3.0150 0.1425 3.0750 0.2025 ;
        RECT 3.0150 0.8325 3.0750 0.8925 ;
        RECT 2.9100 0.4875 2.9700 0.5475 ;
        RECT 2.8050 0.1575 2.8650 0.2175 ;
        RECT 2.8050 0.6675 2.8650 0.7275 ;
        RECT 2.7000 0.4875 2.7600 0.5475 ;
        RECT 2.5950 0.1425 2.6550 0.2025 ;
        RECT 2.5950 0.8325 2.6550 0.8925 ;
        RECT 2.4900 0.4875 2.5500 0.5475 ;
        RECT 2.3850 0.1575 2.4450 0.2175 ;
        RECT 2.3850 0.6675 2.4450 0.7275 ;
        RECT 2.2800 0.4875 2.3400 0.5475 ;
        RECT 2.1750 0.1425 2.2350 0.2025 ;
        RECT 2.1750 0.8325 2.2350 0.8925 ;
        RECT 2.0700 0.4875 2.1300 0.5475 ;
        RECT 1.9650 0.1575 2.0250 0.2175 ;
        RECT 1.9650 0.6675 2.0250 0.7275 ;
        RECT 1.8600 0.4875 1.9200 0.5475 ;
        RECT 1.7550 0.1425 1.8150 0.2025 ;
        RECT 1.7550 0.8325 1.8150 0.8925 ;
        RECT 1.6500 0.4875 1.7100 0.5475 ;
        RECT 1.5450 0.1575 1.6050 0.2175 ;
        RECT 1.5450 0.6675 1.6050 0.7275 ;
        RECT 1.4400 0.4875 1.5000 0.5475 ;
        RECT 1.3350 0.1425 1.3950 0.2025 ;
        RECT 1.3350 0.8325 1.3950 0.8925 ;
        RECT 1.2300 0.4875 1.2900 0.5475 ;
        RECT 1.1250 0.1575 1.1850 0.2175 ;
        RECT 1.1250 0.6675 1.1850 0.7275 ;
        RECT 1.0200 0.4875 1.0800 0.5475 ;
        RECT 0.9150 0.1425 0.9750 0.2025 ;
        RECT 0.9150 0.8325 0.9750 0.8925 ;
        RECT 0.8100 0.4875 0.8700 0.5475 ;
        RECT 0.7050 0.1575 0.7650 0.2175 ;
        RECT 0.7050 0.6675 0.7650 0.7275 ;
        RECT 0.6000 0.4875 0.6600 0.5475 ;
        RECT 0.4950 0.1425 0.5550 0.2025 ;
        RECT 0.4950 0.8325 0.5550 0.8925 ;
        RECT 0.3900 0.4875 0.4500 0.5475 ;
        RECT 0.2850 0.1575 0.3450 0.2175 ;
        RECT 0.2850 0.6675 0.3450 0.7275 ;
        RECT 0.1800 0.4875 0.2400 0.5475 ;
        RECT 0.0750 0.1575 0.1350 0.2175 ;
        RECT 0.0750 0.8025 0.1350 0.8625 ;
        LAYER M1 ;
        RECT 10.3575 0.6675 10.4325 0.8250 ;
        RECT 7.0800 0.4650 10.3650 0.5700 ;
        RECT 3.6000 0.6675 10.3575 0.7425 ;
        RECT 10.1325 0.1500 10.2375 0.3900 ;
        RECT 9.8175 0.2925 10.1325 0.3900 ;
        RECT 9.7125 0.1500 9.8175 0.3900 ;
        RECT 9.3975 0.2925 9.7125 0.3900 ;
        RECT 9.2925 0.1500 9.3975 0.3900 ;
        RECT 8.9775 0.2925 9.2925 0.3900 ;
        RECT 8.8725 0.1500 8.9775 0.3900 ;
        RECT 8.5575 0.2925 8.8725 0.3900 ;
        RECT 8.4525 0.1500 8.5575 0.3900 ;
        RECT 8.1450 0.2925 8.4525 0.3900 ;
        RECT 8.0250 0.1500 8.1450 0.3900 ;
        RECT 7.7250 0.2925 8.0250 0.3900 ;
        RECT 7.6050 0.1500 7.7250 0.3900 ;
        RECT 7.3050 0.2925 7.6050 0.3900 ;
        RECT 7.1850 0.1500 7.3050 0.3900 ;
        RECT 6.6750 0.2925 7.1850 0.3900 ;
        RECT 0.1575 0.8250 6.9000 0.9000 ;
        RECT 3.5175 0.4650 6.8100 0.5700 ;
        RECT 6.5550 0.1500 6.6750 0.3900 ;
        RECT 6.2550 0.2925 6.5550 0.3900 ;
        RECT 6.1350 0.1500 6.2550 0.3900 ;
        RECT 5.8350 0.2925 6.1350 0.3900 ;
        RECT 5.7150 0.1500 5.8350 0.3900 ;
        RECT 5.4150 0.2925 5.7150 0.3900 ;
        RECT 5.2950 0.1500 5.4150 0.3900 ;
        RECT 4.9950 0.2925 5.2950 0.3900 ;
        RECT 4.8750 0.1500 4.9950 0.3900 ;
        RECT 4.5750 0.2925 4.8750 0.3900 ;
        RECT 4.4550 0.1500 4.5750 0.3900 ;
        RECT 4.1550 0.2925 4.4550 0.3900 ;
        RECT 4.0350 0.1500 4.1550 0.3900 ;
        RECT 3.7350 0.2925 4.0350 0.3900 ;
        RECT 3.6150 0.1500 3.7350 0.3900 ;
        RECT 3.3150 0.2925 3.6150 0.3900 ;
        RECT 3.1950 0.1500 3.3150 0.3900 ;
        RECT 0.2625 0.6450 3.3150 0.7500 ;
        RECT 2.8950 0.2925 3.1950 0.3900 ;
        RECT 2.7750 0.1500 2.8950 0.3900 ;
        RECT 2.4750 0.2925 2.7750 0.3900 ;
        RECT 2.3550 0.1500 2.4750 0.3900 ;
        RECT 2.0550 0.2925 2.3550 0.3900 ;
        RECT 1.9350 0.1500 2.0550 0.3900 ;
        RECT 1.6350 0.2925 1.9350 0.3900 ;
        RECT 1.5150 0.1500 1.6350 0.3900 ;
        RECT 1.2150 0.2925 1.5150 0.3900 ;
        RECT 1.0950 0.1500 1.2150 0.3900 ;
        RECT 0.7950 0.2925 1.0950 0.3900 ;
        RECT 0.6750 0.1500 0.7950 0.3900 ;
        RECT 0.3750 0.2925 0.6750 0.3900 ;
        RECT 0.2550 0.1500 0.3750 0.3900 ;
        RECT 0.0525 0.7725 0.1575 0.9000 ;
        LAYER M2 ;
        RECT 1.9725 0.2775 2.1000 0.3975 ;
        RECT 1.9725 0.6375 2.1000 0.7575 ;
        RECT 1.4700 0.2775 1.5975 0.3975 ;
        RECT 1.4700 0.6375 1.5975 0.7575 ;
    END
END NR3_0100


MACRO NR3_0111
    CLASS CORE ;
    FOREIGN NR3_0111 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.4600 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 0.7875 0.2625 1.1025 0.7800 ;
        VIA 0.9450 0.3450 VIA12_slot ;
        VIA 0.9450 0.6975 VIA12_slot ;
        END
    END ZN
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 4.5075 0.4125 4.5825 0.5775 ;
        RECT 4.0425 0.4125 4.5075 0.4875 ;
        VIA 4.5450 0.4950 VIA12_square ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 2.5875 0.4125 2.6625 0.5775 ;
        RECT 2.1225 0.4125 2.5875 0.4875 ;
        VIA 2.6250 0.4950 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1425 0.4575 1.7400 0.5625 ;
        RECT 0.0675 0.3675 0.1425 0.6825 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 5.4075 -0.0750 5.4600 0.0750 ;
        RECT 5.3025 -0.0750 5.4075 0.2625 ;
        RECT 4.9950 -0.0750 5.3025 0.0750 ;
        RECT 4.8750 -0.0750 4.9950 0.1950 ;
        RECT 4.5750 -0.0750 4.8750 0.0750 ;
        RECT 4.4550 -0.0750 4.5750 0.1950 ;
        RECT 4.1550 -0.0750 4.4550 0.0750 ;
        RECT 4.0350 -0.0750 4.1550 0.1950 ;
        RECT 3.7350 -0.0750 4.0350 0.0750 ;
        RECT 3.6150 -0.0750 3.7350 0.2175 ;
        RECT 3.5250 -0.0750 3.6150 0.0750 ;
        RECT 3.4050 -0.0750 3.5250 0.2175 ;
        RECT 3.1050 -0.0750 3.4050 0.0750 ;
        RECT 2.9850 -0.0750 3.1050 0.1950 ;
        RECT 2.6850 -0.0750 2.9850 0.0750 ;
        RECT 2.5650 -0.0750 2.6850 0.1950 ;
        RECT 2.2650 -0.0750 2.5650 0.0750 ;
        RECT 2.1450 -0.0750 2.2650 0.1950 ;
        RECT 1.8450 -0.0750 2.1450 0.0750 ;
        RECT 1.7250 -0.0750 1.8450 0.1950 ;
        RECT 1.4250 -0.0750 1.7250 0.0750 ;
        RECT 1.3050 -0.0750 1.4250 0.1950 ;
        RECT 1.0050 -0.0750 1.3050 0.0750 ;
        RECT 0.8850 -0.0750 1.0050 0.1950 ;
        RECT 0.5850 -0.0750 0.8850 0.0750 ;
        RECT 0.4650 -0.0750 0.5850 0.1950 ;
        RECT 0.1650 -0.0750 0.4650 0.0750 ;
        RECT 0.0450 -0.0750 0.1650 0.2250 ;
        RECT 0.0000 -0.0750 0.0450 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 5.2050 0.9750 5.4600 1.1250 ;
        RECT 5.0850 0.8175 5.2050 1.1250 ;
        RECT 4.7850 0.9750 5.0850 1.1250 ;
        RECT 4.6650 0.8175 4.7850 1.1250 ;
        RECT 4.3650 0.9750 4.6650 1.1250 ;
        RECT 4.2450 0.8175 4.3650 1.1250 ;
        RECT 3.9450 0.9750 4.2450 1.1250 ;
        RECT 3.8250 0.8175 3.9450 1.1250 ;
        RECT 0.0000 0.9750 3.8250 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 5.3250 0.1725 5.3850 0.2325 ;
        RECT 5.3250 0.7350 5.3850 0.7950 ;
        RECT 5.2200 0.4875 5.2800 0.5475 ;
        RECT 5.1150 0.2775 5.1750 0.3375 ;
        RECT 5.1150 0.8400 5.1750 0.9000 ;
        RECT 5.0100 0.4875 5.0700 0.5475 ;
        RECT 4.9050 0.1275 4.9650 0.1875 ;
        RECT 4.9050 0.6750 4.9650 0.7350 ;
        RECT 4.8000 0.4875 4.8600 0.5475 ;
        RECT 4.6950 0.3075 4.7550 0.3675 ;
        RECT 4.6950 0.8400 4.7550 0.9000 ;
        RECT 4.5900 0.4875 4.6500 0.5475 ;
        RECT 4.4850 0.1275 4.5450 0.1875 ;
        RECT 4.4850 0.6750 4.5450 0.7350 ;
        RECT 4.3800 0.4875 4.4400 0.5475 ;
        RECT 4.2750 0.3075 4.3350 0.3675 ;
        RECT 4.2750 0.8400 4.3350 0.9000 ;
        RECT 4.1700 0.4875 4.2300 0.5475 ;
        RECT 4.0650 0.1275 4.1250 0.1875 ;
        RECT 4.0650 0.6750 4.1250 0.7350 ;
        RECT 3.9600 0.4875 4.0200 0.5475 ;
        RECT 3.8550 0.3075 3.9150 0.3675 ;
        RECT 3.8550 0.8400 3.9150 0.9000 ;
        RECT 3.7500 0.4875 3.8100 0.5475 ;
        RECT 3.6450 0.1575 3.7050 0.2175 ;
        RECT 3.6450 0.6750 3.7050 0.7350 ;
        RECT 3.4350 0.1575 3.4950 0.2175 ;
        RECT 3.4350 0.8325 3.4950 0.8925 ;
        RECT 3.3300 0.4875 3.3900 0.5475 ;
        RECT 3.2250 0.3075 3.2850 0.3675 ;
        RECT 3.2250 0.6750 3.2850 0.7350 ;
        RECT 3.1200 0.4875 3.1800 0.5475 ;
        RECT 3.0150 0.1275 3.0750 0.1875 ;
        RECT 3.0150 0.8325 3.0750 0.8925 ;
        RECT 2.9100 0.4875 2.9700 0.5475 ;
        RECT 2.8050 0.3075 2.8650 0.3675 ;
        RECT 2.8050 0.6750 2.8650 0.7350 ;
        RECT 2.7000 0.4875 2.7600 0.5475 ;
        RECT 2.5950 0.1275 2.6550 0.1875 ;
        RECT 2.5950 0.8325 2.6550 0.8925 ;
        RECT 2.4900 0.4875 2.5500 0.5475 ;
        RECT 2.3850 0.3075 2.4450 0.3675 ;
        RECT 2.3850 0.6750 2.4450 0.7350 ;
        RECT 2.2800 0.4875 2.3400 0.5475 ;
        RECT 2.1750 0.1275 2.2350 0.1875 ;
        RECT 2.1750 0.8325 2.2350 0.8925 ;
        RECT 2.0700 0.4875 2.1300 0.5475 ;
        RECT 1.9650 0.3075 2.0250 0.3675 ;
        RECT 1.9650 0.6750 2.0250 0.7350 ;
        RECT 1.8600 0.4875 1.9200 0.5475 ;
        RECT 1.7550 0.1275 1.8150 0.1875 ;
        RECT 1.7550 0.8325 1.8150 0.8925 ;
        RECT 1.6500 0.4800 1.7100 0.5400 ;
        RECT 1.5450 0.3075 1.6050 0.3675 ;
        RECT 1.5450 0.6675 1.6050 0.7275 ;
        RECT 1.4400 0.4800 1.5000 0.5400 ;
        RECT 1.3350 0.1275 1.3950 0.1875 ;
        RECT 1.3350 0.8325 1.3950 0.8925 ;
        RECT 1.2300 0.4800 1.2900 0.5400 ;
        RECT 1.1250 0.3075 1.1850 0.3675 ;
        RECT 1.1250 0.6675 1.1850 0.7275 ;
        RECT 1.0200 0.4800 1.0800 0.5400 ;
        RECT 0.9150 0.1275 0.9750 0.1875 ;
        RECT 0.9150 0.8325 0.9750 0.8925 ;
        RECT 0.8100 0.4800 0.8700 0.5400 ;
        RECT 0.7050 0.3075 0.7650 0.3675 ;
        RECT 0.7050 0.6675 0.7650 0.7275 ;
        RECT 0.6000 0.4800 0.6600 0.5400 ;
        RECT 0.4950 0.1275 0.5550 0.1875 ;
        RECT 0.4950 0.8325 0.5550 0.8925 ;
        RECT 0.3900 0.4800 0.4500 0.5400 ;
        RECT 0.2850 0.3075 0.3450 0.3675 ;
        RECT 0.2850 0.6675 0.3450 0.7275 ;
        RECT 0.1800 0.4800 0.2400 0.5400 ;
        RECT 0.0750 0.1575 0.1350 0.2175 ;
        RECT 0.0750 0.8175 0.1350 0.8775 ;
        LAYER M1 ;
        RECT 5.3175 0.6675 5.3925 0.8250 ;
        RECT 1.9200 0.6675 5.3175 0.7425 ;
        RECT 3.7425 0.4575 5.2875 0.5775 ;
        RECT 5.0925 0.2550 5.1975 0.3825 ;
        RECT 0.2550 0.3075 5.0925 0.3825 ;
        RECT 0.1575 0.8250 3.5400 0.9000 ;
        RECT 1.8525 0.4575 3.4050 0.5775 ;
        RECT 0.2625 0.6450 1.6350 0.7500 ;
        RECT 0.0525 0.7950 0.1575 0.9000 ;
    END
END NR3_0111


MACRO NR3_1000
    CLASS CORE ;
    FOREIGN NR3_1000 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.8400 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.7275 0.1500 0.8025 0.9000 ;
        RECT 0.6750 0.1500 0.7275 0.3750 ;
        RECT 0.6975 0.6675 0.7275 0.9000 ;
        RECT 0.6150 0.2550 0.6750 0.3750 ;
        RECT 0.3675 0.2550 0.6150 0.3300 ;
        RECT 0.2625 0.1500 0.3675 0.3300 ;
        END
    END ZN
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1425 0.4500 0.2325 0.6000 ;
        RECT 0.0675 0.3675 0.1425 0.6825 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.3825 0.4125 0.4725 0.5175 ;
        RECT 0.3075 0.4125 0.3825 0.8325 ;
        RECT 0.2775 0.6675 0.3075 0.8325 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.6225 0.4500 0.6525 0.5925 ;
        RECT 0.5475 0.4500 0.6225 0.8325 ;
        RECT 0.4875 0.6675 0.5475 0.8325 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.5850 -0.0750 0.8400 0.0750 ;
        RECT 0.4650 -0.0750 0.5850 0.1800 ;
        RECT 0.1425 -0.0750 0.4650 0.0750 ;
        RECT 0.0675 -0.0750 0.1425 0.2475 ;
        RECT 0.0000 -0.0750 0.0675 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.1425 0.9750 0.8400 1.1250 ;
        RECT 0.0675 0.8025 0.1425 1.1250 ;
        RECT 0.0000 0.9750 0.0675 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 0.7050 0.1575 0.7650 0.2175 ;
        RECT 0.7050 0.7575 0.7650 0.8175 ;
        RECT 0.5925 0.4950 0.6525 0.5550 ;
        RECT 0.4950 0.1200 0.5550 0.1800 ;
        RECT 0.3825 0.4200 0.4425 0.4800 ;
        RECT 0.2850 0.1725 0.3450 0.2325 ;
        RECT 0.1725 0.4950 0.2325 0.5550 ;
        RECT 0.0750 0.1575 0.1350 0.2175 ;
        RECT 0.0750 0.8325 0.1350 0.8925 ;
    END
END NR3_1000


MACRO NR3_1010
    CLASS CORE ;
    FOREIGN NR3_1010 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.4700 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 0.9675 0.7125 1.2075 0.7875 ;
        RECT 0.8925 0.2625 0.9675 0.7875 ;
        RECT 0.6525 0.2625 0.8925 0.3375 ;
        VIA 0.9300 0.6825 VIA12_square ;
        VIA 0.8100 0.3000 VIA12_square ;
        END
    END ZN
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.2300 0.4200 1.3350 0.7200 ;
        RECT 1.2150 0.6450 1.2300 0.7200 ;
        RECT 1.1400 0.6450 1.2150 0.8700 ;
        RECT 0.3225 0.7950 1.1400 0.8700 ;
        RECT 0.2475 0.6450 0.3225 0.8700 ;
        RECT 0.1425 0.6450 0.2475 0.7200 ;
        RECT 0.1425 0.4200 0.2325 0.5550 ;
        RECT 0.0675 0.3675 0.1425 0.7200 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.0425 0.1125 1.1175 0.5775 ;
        RECT 0.5325 0.1125 1.0425 0.1875 ;
        RECT 0.4575 0.1125 0.5325 0.4875 ;
        RECT 0.3075 0.4125 0.4575 0.4875 ;
        VIA 1.0800 0.4650 VIA12_square ;
        VIA 0.4200 0.4500 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.7125 0.4200 0.8175 0.6375 ;
        RECT 0.3525 0.5625 0.7125 0.6375 ;
        VIA 0.7650 0.4950 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.4250 -0.0750 1.4700 0.0750 ;
        RECT 1.3050 -0.0750 1.4250 0.2475 ;
        RECT 1.0050 -0.0750 1.3050 0.0750 ;
        RECT 0.8850 -0.0750 1.0050 0.1875 ;
        RECT 0.5850 -0.0750 0.8850 0.0750 ;
        RECT 0.4650 -0.0750 0.5850 0.1875 ;
        RECT 0.1650 -0.0750 0.4650 0.0750 ;
        RECT 0.0450 -0.0750 0.1650 0.2475 ;
        RECT 0.0000 -0.0750 0.0450 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.4175 0.9750 1.4700 1.1250 ;
        RECT 1.3125 0.8100 1.4175 1.1250 ;
        RECT 0.1575 0.9750 1.3125 1.1250 ;
        RECT 0.0525 0.8100 0.1575 1.1250 ;
        RECT 0.0000 0.9750 0.0525 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.3350 0.1575 1.3950 0.2175 ;
        RECT 1.3350 0.8325 1.3950 0.8925 ;
        RECT 1.2300 0.4650 1.2900 0.5250 ;
        RECT 1.1250 0.1800 1.1850 0.2400 ;
        RECT 1.0200 0.4650 1.0800 0.5250 ;
        RECT 0.9150 0.1275 0.9750 0.1875 ;
        RECT 0.8100 0.4650 0.8700 0.5250 ;
        RECT 0.7050 0.1800 0.7650 0.2400 ;
        RECT 0.7050 0.6525 0.7650 0.7125 ;
        RECT 0.6000 0.4650 0.6600 0.5250 ;
        RECT 0.4950 0.1275 0.5550 0.1875 ;
        RECT 0.3900 0.4650 0.4500 0.5250 ;
        RECT 0.2850 0.1800 0.3450 0.2400 ;
        RECT 0.1725 0.4650 0.2325 0.5250 ;
        RECT 0.0750 0.1575 0.1350 0.2175 ;
        RECT 0.0750 0.8325 0.1350 0.8925 ;
        LAYER M1 ;
        RECT 1.1025 0.1575 1.2075 0.3375 ;
        RECT 0.9450 0.4125 1.1550 0.5700 ;
        RECT 0.7875 0.2625 1.1025 0.3375 ;
        RECT 0.6000 0.6450 1.0200 0.7200 ;
        RECT 0.6000 0.4350 0.8700 0.5550 ;
        RECT 0.6825 0.1575 0.7875 0.3375 ;
        RECT 0.3675 0.2625 0.6825 0.3375 ;
        RECT 0.3075 0.4125 0.5250 0.5700 ;
        RECT 0.2625 0.1575 0.3675 0.3375 ;
    END
END NR3_1010


MACRO NR4_0001
    CLASS CORE ;
    FOREIGN NR4_0001 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.4600 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 5.0925 0.1500 5.1975 0.3825 ;
        RECT 4.7775 0.2925 5.0925 0.3825 ;
        RECT 4.6725 0.1500 4.7775 0.3825 ;
        RECT 4.3575 0.2925 4.6725 0.3825 ;
        RECT 4.2525 0.1500 4.3575 0.3825 ;
        RECT 3.9375 0.2925 4.2525 0.3825 ;
        RECT 3.8325 0.1500 3.9375 0.3825 ;
        RECT 3.5175 0.2925 3.8325 0.3825 ;
        RECT 3.4125 0.1500 3.5175 0.3825 ;
        RECT 3.0975 0.2925 3.4125 0.3825 ;
        RECT 2.9925 0.1500 3.0975 0.3825 ;
        RECT 2.4675 0.2925 2.9925 0.3825 ;
        RECT 2.3625 0.1500 2.4675 0.3825 ;
        RECT 2.0475 0.2925 2.3625 0.3825 ;
        RECT 1.9425 0.1500 2.0475 0.3825 ;
        RECT 1.6275 0.2925 1.9425 0.3825 ;
        RECT 1.5225 0.1500 1.6275 0.3825 ;
        RECT 1.2075 0.2925 1.5225 0.3825 ;
        RECT 0.2625 0.6450 1.2150 0.7500 ;
        RECT 1.1025 0.1500 1.2075 0.3825 ;
        RECT 0.7875 0.2925 1.1025 0.3825 ;
        RECT 0.6825 0.1500 0.7875 0.3825 ;
        RECT 0.6375 0.2925 0.6825 0.3825 ;
        RECT 0.3675 0.2925 0.6375 0.3750 ;
        RECT 0.2625 0.1500 0.3675 0.3750 ;
        RECT 0.1125 0.3000 0.2625 0.3750 ;
        RECT 0.1125 0.6450 0.2625 0.7200 ;
        RECT 0.0375 0.3000 0.1125 0.7200 ;
        END
    END ZN
    PIN A4
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 4.4400 0.4125 4.5450 0.6375 ;
        RECT 3.9750 0.4125 4.4400 0.4875 ;
        VIA 4.4925 0.5100 VIA12_square ;
        END
    END A4
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 3.3075 0.5625 3.7725 0.6375 ;
        RECT 3.2025 0.4125 3.3075 0.6375 ;
        VIA 3.2550 0.5025 VIA12_square ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.8375 0.5625 2.3025 0.6375 ;
        RECT 1.7325 0.4125 1.8375 0.6375 ;
        VIA 1.7850 0.5025 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.6600 0.5625 1.1250 0.6375 ;
        RECT 0.5550 0.4125 0.6600 0.6375 ;
        VIA 0.6075 0.5025 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 5.4075 -0.0750 5.4600 0.0750 ;
        RECT 5.3025 -0.0750 5.4075 0.2625 ;
        RECT 4.9950 -0.0750 5.3025 0.0750 ;
        RECT 4.8750 -0.0750 4.9950 0.2100 ;
        RECT 4.5750 -0.0750 4.8750 0.0750 ;
        RECT 4.4550 -0.0750 4.5750 0.2100 ;
        RECT 4.1550 -0.0750 4.4550 0.0750 ;
        RECT 4.0350 -0.0750 4.1550 0.2100 ;
        RECT 3.7350 -0.0750 4.0350 0.0750 ;
        RECT 3.6150 -0.0750 3.7350 0.2100 ;
        RECT 3.3150 -0.0750 3.6150 0.0750 ;
        RECT 3.1950 -0.0750 3.3150 0.2100 ;
        RECT 2.8950 -0.0750 3.1950 0.0750 ;
        RECT 2.7750 -0.0750 2.8950 0.2175 ;
        RECT 2.6850 -0.0750 2.7750 0.0750 ;
        RECT 2.5650 -0.0750 2.6850 0.2175 ;
        RECT 2.2650 -0.0750 2.5650 0.0750 ;
        RECT 2.1450 -0.0750 2.2650 0.2100 ;
        RECT 1.8450 -0.0750 2.1450 0.0750 ;
        RECT 1.7250 -0.0750 1.8450 0.2100 ;
        RECT 1.4175 -0.0750 1.7250 0.0750 ;
        RECT 1.3125 -0.0750 1.4175 0.2175 ;
        RECT 1.0050 -0.0750 1.3125 0.0750 ;
        RECT 0.8850 -0.0750 1.0050 0.2100 ;
        RECT 0.5775 -0.0750 0.8850 0.0750 ;
        RECT 0.4725 -0.0750 0.5775 0.2175 ;
        RECT 0.1650 -0.0750 0.4725 0.0750 ;
        RECT 0.0450 -0.0750 0.1650 0.2250 ;
        RECT 0.0000 -0.0750 0.0450 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 5.2050 0.9750 5.4600 1.1250 ;
        RECT 5.0850 0.8175 5.2050 1.1250 ;
        RECT 4.7850 0.9750 5.0850 1.1250 ;
        RECT 4.6650 0.8175 4.7850 1.1250 ;
        RECT 4.3650 0.9750 4.6650 1.1250 ;
        RECT 4.2450 0.8175 4.3650 1.1250 ;
        RECT 0.0000 0.9750 4.2450 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 5.3250 0.1575 5.3850 0.2175 ;
        RECT 5.3250 0.7350 5.3850 0.7950 ;
        RECT 5.2200 0.4725 5.2800 0.5325 ;
        RECT 5.1150 0.1725 5.1750 0.2325 ;
        RECT 5.1150 0.8400 5.1750 0.9000 ;
        RECT 5.0100 0.4725 5.0700 0.5325 ;
        RECT 4.9050 0.1425 4.9650 0.2025 ;
        RECT 4.9050 0.6750 4.9650 0.7350 ;
        RECT 4.8000 0.4725 4.8600 0.5325 ;
        RECT 4.6950 0.1725 4.7550 0.2325 ;
        RECT 4.6950 0.8400 4.7550 0.9000 ;
        RECT 4.5900 0.4725 4.6500 0.5325 ;
        RECT 4.4850 0.1425 4.5450 0.2025 ;
        RECT 4.4850 0.6750 4.5450 0.7350 ;
        RECT 4.3800 0.4725 4.4400 0.5325 ;
        RECT 4.2750 0.1725 4.3350 0.2325 ;
        RECT 4.2750 0.8400 4.3350 0.9000 ;
        RECT 4.1700 0.4725 4.2300 0.5325 ;
        RECT 4.0650 0.1425 4.1250 0.2025 ;
        RECT 4.0650 0.6750 4.1250 0.7350 ;
        RECT 3.9600 0.4725 4.0200 0.5325 ;
        RECT 3.8550 0.1725 3.9150 0.2325 ;
        RECT 3.8550 0.8325 3.9150 0.8925 ;
        RECT 3.7500 0.4725 3.8100 0.5325 ;
        RECT 3.6450 0.1425 3.7050 0.2025 ;
        RECT 3.6450 0.6750 3.7050 0.7350 ;
        RECT 3.5400 0.4725 3.6000 0.5325 ;
        RECT 3.4350 0.1725 3.4950 0.2325 ;
        RECT 3.4350 0.8325 3.4950 0.8925 ;
        RECT 3.3300 0.4725 3.3900 0.5325 ;
        RECT 3.2250 0.1425 3.2850 0.2025 ;
        RECT 3.2250 0.6750 3.2850 0.7350 ;
        RECT 3.1200 0.4725 3.1800 0.5325 ;
        RECT 3.0150 0.1725 3.0750 0.2325 ;
        RECT 3.0150 0.8325 3.0750 0.8925 ;
        RECT 2.9100 0.4725 2.9700 0.5325 ;
        RECT 2.8050 0.1575 2.8650 0.2175 ;
        RECT 2.8050 0.6600 2.8650 0.7200 ;
        RECT 2.5950 0.1575 2.6550 0.2175 ;
        RECT 2.5950 0.6600 2.6550 0.7200 ;
        RECT 2.4900 0.4800 2.5500 0.5400 ;
        RECT 2.3850 0.1725 2.4450 0.2325 ;
        RECT 2.3850 0.8325 2.4450 0.8925 ;
        RECT 2.2800 0.4800 2.3400 0.5400 ;
        RECT 2.1750 0.1425 2.2350 0.2025 ;
        RECT 2.1750 0.6750 2.2350 0.7350 ;
        RECT 2.0700 0.4800 2.1300 0.5400 ;
        RECT 1.9650 0.1725 2.0250 0.2325 ;
        RECT 1.9650 0.8325 2.0250 0.8925 ;
        RECT 1.8600 0.4800 1.9200 0.5400 ;
        RECT 1.7550 0.1425 1.8150 0.2025 ;
        RECT 1.7550 0.6750 1.8150 0.7350 ;
        RECT 1.6500 0.4800 1.7100 0.5400 ;
        RECT 1.5450 0.1725 1.6050 0.2325 ;
        RECT 1.5450 0.8325 1.6050 0.8925 ;
        RECT 1.4400 0.4800 1.5000 0.5400 ;
        RECT 1.3350 0.1350 1.3950 0.1950 ;
        RECT 1.3350 0.7575 1.3950 0.8175 ;
        RECT 1.2300 0.4800 1.2900 0.5400 ;
        RECT 1.1250 0.1725 1.1850 0.2325 ;
        RECT 1.1250 0.6675 1.1850 0.7275 ;
        RECT 1.0200 0.4725 1.0800 0.5325 ;
        RECT 0.9150 0.1425 0.9750 0.2025 ;
        RECT 0.9150 0.8325 0.9750 0.8925 ;
        RECT 0.8100 0.4800 0.8700 0.5400 ;
        RECT 0.7050 0.1725 0.7650 0.2325 ;
        RECT 0.7050 0.6675 0.7650 0.7275 ;
        RECT 0.6000 0.4725 0.6600 0.5325 ;
        RECT 0.4950 0.1350 0.5550 0.1950 ;
        RECT 0.4950 0.8325 0.5550 0.8925 ;
        RECT 0.3900 0.4725 0.4500 0.5325 ;
        RECT 0.2850 0.1725 0.3450 0.2325 ;
        RECT 0.2850 0.6675 0.3450 0.7275 ;
        RECT 0.1875 0.4800 0.2475 0.5400 ;
        RECT 0.0750 0.1575 0.1350 0.2175 ;
        RECT 0.0750 0.8175 0.1350 0.8775 ;
        LAYER M1 ;
        RECT 5.3175 0.6675 5.3925 0.8250 ;
        RECT 4.1400 0.4575 5.3175 0.5625 ;
        RECT 2.8950 0.6675 5.3175 0.7425 ;
        RECT 2.8800 0.4575 4.0500 0.5625 ;
        RECT 1.5075 0.8250 3.9825 0.9000 ;
        RECT 2.7825 0.6375 2.8950 0.7425 ;
        RECT 2.5725 0.6375 2.6775 0.7425 ;
        RECT 1.4175 0.4575 2.5725 0.5625 ;
        RECT 1.4025 0.6675 2.5725 0.7425 ;
        RECT 1.3275 0.6675 1.4025 0.9000 ;
        RECT 0.1650 0.8250 1.3275 0.9000 ;
        RECT 0.4800 0.4575 1.3125 0.5700 ;
        RECT 0.1875 0.4500 0.4800 0.5700 ;
        RECT 0.0450 0.7950 0.1650 0.9000 ;
    END
END NR4_0001


MACRO NR4_0011
    CLASS CORE ;
    FOREIGN NR4_0011 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.7800 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 3.4125 0.1500 3.5175 0.3825 ;
        RECT 3.0975 0.2925 3.4125 0.3825 ;
        RECT 2.9925 0.1500 3.0975 0.3825 ;
        RECT 2.6775 0.2925 2.9925 0.3825 ;
        RECT 2.5725 0.1500 2.6775 0.3825 ;
        RECT 2.2575 0.2925 2.5725 0.3825 ;
        RECT 2.1525 0.1500 2.2575 0.3825 ;
        RECT 1.6275 0.2925 2.1525 0.3825 ;
        RECT 1.5225 0.1500 1.6275 0.3825 ;
        RECT 1.2075 0.2925 1.5225 0.3825 ;
        RECT 1.1025 0.1500 1.2075 0.3825 ;
        RECT 0.7875 0.2925 1.1025 0.3825 ;
        RECT 0.2625 0.6450 0.7950 0.7500 ;
        RECT 0.6825 0.1500 0.7875 0.3825 ;
        RECT 0.6375 0.2925 0.6825 0.3825 ;
        RECT 0.3675 0.2925 0.6375 0.3750 ;
        RECT 0.2625 0.1500 0.3675 0.3750 ;
        RECT 0.1125 0.3000 0.2625 0.3750 ;
        RECT 0.1125 0.6450 0.2625 0.7200 ;
        RECT 0.0375 0.3000 0.1125 0.7200 ;
        END
    END ZN
    PIN A4
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 3.1800 0.4125 3.2850 0.6375 ;
        RECT 2.7150 0.4125 3.1800 0.4875 ;
        VIA 3.2325 0.5100 VIA12_square ;
        END
    END A4
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 2.4675 0.5625 2.9325 0.6375 ;
        RECT 2.3625 0.4125 2.4675 0.6375 ;
        VIA 2.4150 0.5025 VIA12_square ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.4175 0.5625 1.8825 0.6375 ;
        RECT 1.3125 0.4125 1.4175 0.6375 ;
        VIA 1.3650 0.5025 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.6600 0.5625 1.1250 0.6375 ;
        RECT 0.5550 0.4125 0.6600 0.6375 ;
        VIA 0.6075 0.5025 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 3.7275 -0.0750 3.7800 0.0750 ;
        RECT 3.6225 -0.0750 3.7275 0.2625 ;
        RECT 3.3150 -0.0750 3.6225 0.0750 ;
        RECT 3.1950 -0.0750 3.3150 0.2100 ;
        RECT 2.8950 -0.0750 3.1950 0.0750 ;
        RECT 2.7750 -0.0750 2.8950 0.2100 ;
        RECT 2.4750 -0.0750 2.7750 0.0750 ;
        RECT 2.3550 -0.0750 2.4750 0.2100 ;
        RECT 2.0550 -0.0750 2.3550 0.0750 ;
        RECT 1.9350 -0.0750 2.0550 0.2175 ;
        RECT 1.8450 -0.0750 1.9350 0.0750 ;
        RECT 1.7250 -0.0750 1.8450 0.2175 ;
        RECT 1.4250 -0.0750 1.7250 0.0750 ;
        RECT 1.3050 -0.0750 1.4250 0.2100 ;
        RECT 0.9975 -0.0750 1.3050 0.0750 ;
        RECT 0.8925 -0.0750 0.9975 0.2175 ;
        RECT 0.5775 -0.0750 0.8925 0.0750 ;
        RECT 0.4725 -0.0750 0.5775 0.2175 ;
        RECT 0.1650 -0.0750 0.4725 0.0750 ;
        RECT 0.0450 -0.0750 0.1650 0.2250 ;
        RECT 0.0000 -0.0750 0.0450 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 3.5250 0.9750 3.7800 1.1250 ;
        RECT 3.4050 0.8175 3.5250 1.1250 ;
        RECT 3.1050 0.9750 3.4050 1.1250 ;
        RECT 2.9850 0.8175 3.1050 1.1250 ;
        RECT 0.0000 0.9750 2.9850 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 3.6450 0.1575 3.7050 0.2175 ;
        RECT 3.6450 0.7350 3.7050 0.7950 ;
        RECT 3.5400 0.4725 3.6000 0.5325 ;
        RECT 3.4350 0.1725 3.4950 0.2325 ;
        RECT 3.4350 0.8400 3.4950 0.9000 ;
        RECT 3.3300 0.4725 3.3900 0.5325 ;
        RECT 3.2250 0.1425 3.2850 0.2025 ;
        RECT 3.2250 0.6750 3.2850 0.7350 ;
        RECT 3.1200 0.4725 3.1800 0.5325 ;
        RECT 3.0150 0.1725 3.0750 0.2325 ;
        RECT 3.0150 0.8400 3.0750 0.9000 ;
        RECT 2.9100 0.4725 2.9700 0.5325 ;
        RECT 2.8050 0.1425 2.8650 0.2025 ;
        RECT 2.8050 0.6750 2.8650 0.7350 ;
        RECT 2.7000 0.4725 2.7600 0.5325 ;
        RECT 2.5950 0.1725 2.6550 0.2325 ;
        RECT 2.5950 0.8325 2.6550 0.8925 ;
        RECT 2.4900 0.4725 2.5500 0.5325 ;
        RECT 2.3850 0.1425 2.4450 0.2025 ;
        RECT 2.3850 0.6750 2.4450 0.7350 ;
        RECT 2.2800 0.4725 2.3400 0.5325 ;
        RECT 2.1750 0.1725 2.2350 0.2325 ;
        RECT 2.1750 0.8325 2.2350 0.8925 ;
        RECT 2.0700 0.4725 2.1300 0.5325 ;
        RECT 1.9650 0.1575 2.0250 0.2175 ;
        RECT 1.9650 0.6600 2.0250 0.7200 ;
        RECT 1.7550 0.1575 1.8150 0.2175 ;
        RECT 1.7550 0.6600 1.8150 0.7200 ;
        RECT 1.6500 0.4800 1.7100 0.5400 ;
        RECT 1.5450 0.1725 1.6050 0.2325 ;
        RECT 1.5450 0.8325 1.6050 0.8925 ;
        RECT 1.4400 0.4800 1.5000 0.5400 ;
        RECT 1.3350 0.1425 1.3950 0.2025 ;
        RECT 1.3350 0.6750 1.3950 0.7350 ;
        RECT 1.2300 0.4800 1.2900 0.5400 ;
        RECT 1.1250 0.1725 1.1850 0.2325 ;
        RECT 1.1250 0.8325 1.1850 0.8925 ;
        RECT 1.0200 0.4800 1.0800 0.5400 ;
        RECT 0.9150 0.1350 0.9750 0.1950 ;
        RECT 0.9150 0.7575 0.9750 0.8175 ;
        RECT 0.8100 0.4800 0.8700 0.5400 ;
        RECT 0.7050 0.1725 0.7650 0.2325 ;
        RECT 0.7050 0.6675 0.7650 0.7275 ;
        RECT 0.6000 0.4725 0.6600 0.5325 ;
        RECT 0.4950 0.1350 0.5550 0.1950 ;
        RECT 0.4950 0.8325 0.5550 0.8925 ;
        RECT 0.3900 0.4725 0.4500 0.5325 ;
        RECT 0.2850 0.1725 0.3450 0.2325 ;
        RECT 0.2850 0.6675 0.3450 0.7275 ;
        RECT 0.1875 0.4800 0.2475 0.5400 ;
        RECT 0.0750 0.1575 0.1350 0.2175 ;
        RECT 0.0750 0.8175 0.1350 0.8775 ;
        LAYER M1 ;
        RECT 3.6375 0.6675 3.7125 0.8250 ;
        RECT 2.8800 0.4575 3.6375 0.5625 ;
        RECT 2.0550 0.6675 3.6375 0.7425 ;
        RECT 2.0400 0.4575 2.7900 0.5625 ;
        RECT 1.0875 0.8250 2.7225 0.9000 ;
        RECT 1.9425 0.6375 2.0550 0.7425 ;
        RECT 1.7325 0.6375 1.8375 0.7425 ;
        RECT 0.9975 0.4575 1.7325 0.5625 ;
        RECT 0.9825 0.6675 1.7325 0.7425 ;
        RECT 0.9075 0.6675 0.9825 0.9000 ;
        RECT 0.1650 0.8250 0.9075 0.9000 ;
        RECT 0.4800 0.4575 0.8925 0.5700 ;
        RECT 0.1875 0.4500 0.4800 0.5700 ;
        RECT 0.0450 0.7950 0.1650 0.9000 ;
    END
END NR4_0011


MACRO NR4_0100
    CLASS CORE ;
    FOREIGN NR4_0100 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.3600 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 1.9425 0.2625 2.1000 0.3825 ;
        RECT 1.9425 0.6600 2.1000 0.7800 ;
        RECT 1.6275 0.2625 1.9425 0.7800 ;
        RECT 1.4700 0.2625 1.6275 0.3825 ;
        RECT 1.4700 0.6600 1.6275 0.7800 ;
        VIA 1.9425 0.3225 VIA12_slot ;
        VIA 1.9425 0.7200 VIA12_slot ;
        VIA 1.6275 0.3225 VIA12_slot ;
        VIA 1.6275 0.7200 VIA12_slot ;
        END
    END ZN
    PIN A4
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.7050 0.4125 1.1700 0.4875 ;
        VIA 0.8625 0.4500 VIA12_square ;
        END
    END A4
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.5550 0.5625 1.0200 0.6375 ;
        VIA 0.6675 0.6000 VIA12_square ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.3525 0.7125 0.8175 0.7875 ;
        VIA 0.4650 0.7500 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.4275 0.1125 0.9450 0.1875 ;
        RECT 0.3525 0.1125 0.4275 0.6375 ;
        RECT 0.1575 0.5625 0.3525 0.6375 ;
        VIA 0.2550 0.6000 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 3.1050 -0.0750 3.3600 0.0750 ;
        RECT 2.9850 -0.0750 3.1050 0.1875 ;
        RECT 2.6850 -0.0750 2.9850 0.0750 ;
        RECT 2.5650 -0.0750 2.6850 0.1875 ;
        RECT 2.2650 -0.0750 2.5650 0.0750 ;
        RECT 2.1450 -0.0750 2.2650 0.1875 ;
        RECT 1.8450 -0.0750 2.1450 0.0750 ;
        RECT 1.7250 -0.0750 1.8450 0.1875 ;
        RECT 1.4250 -0.0750 1.7250 0.0750 ;
        RECT 1.3050 -0.0750 1.4250 0.1875 ;
        RECT 0.9825 -0.0750 1.3050 0.0750 ;
        RECT 0.9075 -0.0750 0.9825 0.2475 ;
        RECT 0.5850 -0.0750 0.9075 0.0750 ;
        RECT 0.4650 -0.0750 0.5850 0.1800 ;
        RECT 0.1650 -0.0750 0.4650 0.0750 ;
        RECT 0.0450 -0.0750 0.1650 0.2175 ;
        RECT 0.0000 -0.0750 0.0450 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 3.0975 0.9750 3.3600 1.1250 ;
        RECT 2.9925 0.8100 3.0975 1.1250 ;
        RECT 2.6850 0.9750 2.9925 1.1250 ;
        RECT 2.5650 0.8175 2.6850 1.1250 ;
        RECT 2.2650 0.9750 2.5650 1.1250 ;
        RECT 2.1450 0.8550 2.2650 1.1250 ;
        RECT 1.8450 0.9750 2.1450 1.1250 ;
        RECT 1.7250 0.8550 1.8450 1.1250 ;
        RECT 1.4250 0.9750 1.7250 1.1250 ;
        RECT 1.3050 0.8550 1.4250 1.1250 ;
        RECT 0.9825 0.9750 1.3050 1.1250 ;
        RECT 0.9075 0.8025 0.9825 1.1250 ;
        RECT 0.0000 0.9750 0.9075 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 3.2250 0.2250 3.2850 0.2850 ;
        RECT 3.2250 0.7575 3.2850 0.8175 ;
        RECT 3.1200 0.4650 3.1800 0.5250 ;
        RECT 3.0150 0.1275 3.0750 0.1875 ;
        RECT 3.0150 0.8325 3.0750 0.8925 ;
        RECT 2.9100 0.4650 2.9700 0.5250 ;
        RECT 2.8050 0.2700 2.8650 0.3300 ;
        RECT 2.8050 0.6675 2.8650 0.7275 ;
        RECT 2.7000 0.4650 2.7600 0.5250 ;
        RECT 2.5950 0.1275 2.6550 0.1875 ;
        RECT 2.5950 0.8250 2.6550 0.8850 ;
        RECT 2.4900 0.4650 2.5500 0.5250 ;
        RECT 2.3850 0.2850 2.4450 0.3450 ;
        RECT 2.3850 0.6900 2.4450 0.7500 ;
        RECT 2.2800 0.4650 2.3400 0.5250 ;
        RECT 2.1750 0.1275 2.2350 0.1875 ;
        RECT 2.1750 0.8625 2.2350 0.9225 ;
        RECT 2.0700 0.4650 2.1300 0.5250 ;
        RECT 1.9650 0.2850 2.0250 0.3450 ;
        RECT 1.9650 0.6900 2.0250 0.7500 ;
        RECT 1.8600 0.4650 1.9200 0.5250 ;
        RECT 1.7550 0.1275 1.8150 0.1875 ;
        RECT 1.7550 0.8625 1.8150 0.9225 ;
        RECT 1.6500 0.4650 1.7100 0.5250 ;
        RECT 1.5450 0.2850 1.6050 0.3450 ;
        RECT 1.5450 0.6900 1.6050 0.7500 ;
        RECT 1.4400 0.4650 1.5000 0.5250 ;
        RECT 1.3350 0.1275 1.3950 0.1875 ;
        RECT 1.3350 0.8625 1.3950 0.9225 ;
        RECT 1.2300 0.4650 1.2900 0.5250 ;
        RECT 1.1250 0.2850 1.1850 0.3450 ;
        RECT 1.1250 0.6900 1.1850 0.7500 ;
        RECT 1.0200 0.4875 1.0800 0.5475 ;
        RECT 0.9150 0.1575 0.9750 0.2175 ;
        RECT 0.9150 0.8325 0.9750 0.8925 ;
        RECT 0.8175 0.4950 0.8775 0.5550 ;
        RECT 0.7050 0.1725 0.7650 0.2325 ;
        RECT 0.6075 0.4800 0.6675 0.5400 ;
        RECT 0.4950 0.1200 0.5550 0.1800 ;
        RECT 0.3975 0.4950 0.4575 0.5550 ;
        RECT 0.2850 0.1725 0.3450 0.2325 ;
        RECT 0.1875 0.4950 0.2475 0.5550 ;
        RECT 0.0750 0.1575 0.1350 0.2175 ;
        RECT 0.0750 0.7575 0.1350 0.8175 ;
        LAYER M1 ;
        RECT 3.2025 0.1950 3.3075 0.3375 ;
        RECT 3.2175 0.6600 3.2925 0.8700 ;
        RECT 2.8050 0.4125 3.2475 0.5325 ;
        RECT 2.6175 0.6600 3.2175 0.7350 ;
        RECT 2.6175 0.2625 3.2025 0.3375 ;
        RECT 2.7000 0.4125 2.8050 0.5625 ;
        RECT 2.5425 0.2625 2.6175 0.7350 ;
        RECT 1.1250 0.4575 2.5425 0.5325 ;
        RECT 1.1025 0.2625 2.4675 0.3825 ;
        RECT 1.1025 0.6600 2.4675 0.7800 ;
        RECT 1.0200 0.4575 1.1250 0.5850 ;
        RECT 0.7800 0.4125 0.9450 0.6825 ;
        RECT 0.6825 0.1500 0.7875 0.3375 ;
        RECT 0.5775 0.4125 0.7050 0.7275 ;
        RECT 0.3750 0.2550 0.6825 0.3375 ;
        RECT 0.3975 0.4575 0.5025 0.8550 ;
        RECT 0.2625 0.1500 0.3750 0.3825 ;
        RECT 0.2175 0.4575 0.3225 0.7425 ;
        RECT 0.1125 0.3075 0.2625 0.3825 ;
        RECT 0.1875 0.4575 0.2175 0.5925 ;
        RECT 0.1125 0.6675 0.1425 0.9000 ;
        RECT 0.0375 0.3075 0.1125 0.9000 ;
        LAYER VIA1 ;
        RECT 2.7975 0.4125 2.8725 0.4875 ;
        RECT 0.6375 0.2625 0.7125 0.3375 ;
        LAYER M2 ;
        RECT 1.9725 0.2625 2.1000 0.3825 ;
        RECT 1.9725 0.6600 2.1000 0.7800 ;
        RECT 1.4700 0.2625 1.5975 0.3825 ;
        RECT 1.4700 0.6600 1.5975 0.7800 ;
        RECT 2.3250 0.4125 3.0075 0.4875 ;
        RECT 2.2500 0.1125 2.3250 0.4875 ;
        RECT 1.2675 0.1125 2.2500 0.1875 ;
        RECT 1.1925 0.1125 1.2675 0.3375 ;
        RECT 0.5925 0.2625 1.1925 0.3375 ;
    END
END NR4_0100


MACRO NR4_0111
    CLASS CORE ;
    FOREIGN NR4_0111 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.1400 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 0.7875 0.2625 1.1025 0.7800 ;
        VIA 0.9450 0.3450 VIA12_slot ;
        VIA 0.9450 0.6975 VIA12_slot ;
        END
    END ZN
    PIN A4
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 6.3750 0.4125 6.4500 0.5775 ;
        RECT 5.9100 0.4125 6.3750 0.4875 ;
        VIA 6.4125 0.4950 VIA12_square ;
        END
    END A4
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 4.2675 0.4125 4.3425 0.5775 ;
        RECT 3.8025 0.4125 4.2675 0.4875 ;
        VIA 4.3050 0.4950 VIA12_square ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 2.5875 0.4125 2.6625 0.5775 ;
        RECT 2.1225 0.4125 2.5875 0.4875 ;
        VIA 2.6250 0.4950 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1425 0.4650 1.7400 0.5700 ;
        RECT 0.0675 0.3675 0.1425 0.6825 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 7.0875 -0.0750 7.1400 0.0750 ;
        RECT 6.9825 -0.0750 7.0875 0.2625 ;
        RECT 6.6750 -0.0750 6.9825 0.0750 ;
        RECT 6.5550 -0.0750 6.6750 0.2100 ;
        RECT 6.2550 -0.0750 6.5550 0.0750 ;
        RECT 6.1350 -0.0750 6.2550 0.2100 ;
        RECT 5.8350 -0.0750 6.1350 0.0750 ;
        RECT 5.7150 -0.0750 5.8350 0.2100 ;
        RECT 5.4150 -0.0750 5.7150 0.0750 ;
        RECT 5.2950 -0.0750 5.4150 0.2100 ;
        RECT 4.9950 -0.0750 5.2950 0.0750 ;
        RECT 4.8750 -0.0750 4.9950 0.2100 ;
        RECT 4.5750 -0.0750 4.8750 0.0750 ;
        RECT 4.4550 -0.0750 4.5750 0.2100 ;
        RECT 4.1550 -0.0750 4.4550 0.0750 ;
        RECT 4.0350 -0.0750 4.1550 0.2100 ;
        RECT 3.7350 -0.0750 4.0350 0.0750 ;
        RECT 3.6150 -0.0750 3.7350 0.2175 ;
        RECT 3.5250 -0.0750 3.6150 0.0750 ;
        RECT 3.4050 -0.0750 3.5250 0.2175 ;
        RECT 3.1050 -0.0750 3.4050 0.0750 ;
        RECT 2.9850 -0.0750 3.1050 0.1950 ;
        RECT 2.6850 -0.0750 2.9850 0.0750 ;
        RECT 2.5650 -0.0750 2.6850 0.2100 ;
        RECT 2.2650 -0.0750 2.5650 0.0750 ;
        RECT 2.1450 -0.0750 2.2650 0.2100 ;
        RECT 1.8450 -0.0750 2.1450 0.0750 ;
        RECT 1.7250 -0.0750 1.8450 0.2100 ;
        RECT 1.4250 -0.0750 1.7250 0.0750 ;
        RECT 1.3050 -0.0750 1.4250 0.2100 ;
        RECT 1.0050 -0.0750 1.3050 0.0750 ;
        RECT 0.8850 -0.0750 1.0050 0.2100 ;
        RECT 0.5850 -0.0750 0.8850 0.0750 ;
        RECT 0.4650 -0.0750 0.5850 0.2100 ;
        RECT 0.1650 -0.0750 0.4650 0.0750 ;
        RECT 0.0450 -0.0750 0.1650 0.2325 ;
        RECT 0.0000 -0.0750 0.0450 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 6.8850 0.9750 7.1400 1.1250 ;
        RECT 6.7650 0.8175 6.8850 1.1250 ;
        RECT 6.4650 0.9750 6.7650 1.1250 ;
        RECT 6.3450 0.8175 6.4650 1.1250 ;
        RECT 6.0450 0.9750 6.3450 1.1250 ;
        RECT 5.9250 0.8175 6.0450 1.1250 ;
        RECT 5.6250 0.9750 5.9250 1.1250 ;
        RECT 5.5050 0.8175 5.6250 1.1250 ;
        RECT 0.0000 0.9750 5.5050 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 7.0050 0.1725 7.0650 0.2325 ;
        RECT 7.0050 0.7350 7.0650 0.7950 ;
        RECT 6.9000 0.4875 6.9600 0.5475 ;
        RECT 6.7950 0.2775 6.8550 0.3375 ;
        RECT 6.7950 0.8400 6.8550 0.9000 ;
        RECT 6.6900 0.4875 6.7500 0.5475 ;
        RECT 6.5850 0.1425 6.6450 0.2025 ;
        RECT 6.5850 0.6750 6.6450 0.7350 ;
        RECT 6.4800 0.4875 6.5400 0.5475 ;
        RECT 6.3750 0.3075 6.4350 0.3675 ;
        RECT 6.3750 0.8400 6.4350 0.9000 ;
        RECT 6.2700 0.4875 6.3300 0.5475 ;
        RECT 6.1650 0.1425 6.2250 0.2025 ;
        RECT 6.1650 0.6750 6.2250 0.7350 ;
        RECT 6.0600 0.4875 6.1200 0.5475 ;
        RECT 5.9550 0.3075 6.0150 0.3675 ;
        RECT 5.9550 0.8400 6.0150 0.9000 ;
        RECT 5.8500 0.4875 5.9100 0.5475 ;
        RECT 5.7450 0.1425 5.8050 0.2025 ;
        RECT 5.7450 0.6750 5.8050 0.7350 ;
        RECT 5.6400 0.4875 5.7000 0.5475 ;
        RECT 5.5350 0.3075 5.5950 0.3675 ;
        RECT 5.5350 0.8400 5.5950 0.9000 ;
        RECT 5.4300 0.4875 5.4900 0.5475 ;
        RECT 5.3250 0.1425 5.3850 0.2025 ;
        RECT 5.3250 0.6750 5.3850 0.7350 ;
        RECT 5.2200 0.4875 5.2800 0.5475 ;
        RECT 5.1150 0.3075 5.1750 0.3675 ;
        RECT 5.1150 0.8325 5.1750 0.8925 ;
        RECT 5.0100 0.4875 5.0700 0.5475 ;
        RECT 4.9050 0.1425 4.9650 0.2025 ;
        RECT 4.9050 0.6750 4.9650 0.7350 ;
        RECT 4.8000 0.4875 4.8600 0.5475 ;
        RECT 4.6950 0.3075 4.7550 0.3675 ;
        RECT 4.6950 0.8325 4.7550 0.8925 ;
        RECT 4.5900 0.4875 4.6500 0.5475 ;
        RECT 4.4850 0.1425 4.5450 0.2025 ;
        RECT 4.4850 0.6750 4.5450 0.7350 ;
        RECT 4.3800 0.4875 4.4400 0.5475 ;
        RECT 4.2750 0.3075 4.3350 0.3675 ;
        RECT 4.2750 0.8325 4.3350 0.8925 ;
        RECT 4.1700 0.4875 4.2300 0.5475 ;
        RECT 4.0650 0.1425 4.1250 0.2025 ;
        RECT 4.0650 0.6750 4.1250 0.7350 ;
        RECT 3.9600 0.4875 4.0200 0.5475 ;
        RECT 3.8550 0.3075 3.9150 0.3675 ;
        RECT 3.8550 0.8325 3.9150 0.8925 ;
        RECT 3.7500 0.4875 3.8100 0.5475 ;
        RECT 3.6450 0.1575 3.7050 0.2175 ;
        RECT 3.6450 0.6750 3.7050 0.7350 ;
        RECT 3.4350 0.1575 3.4950 0.2175 ;
        RECT 3.4350 0.6825 3.4950 0.7425 ;
        RECT 3.3300 0.4875 3.3900 0.5475 ;
        RECT 3.2250 0.3075 3.2850 0.3675 ;
        RECT 3.2250 0.8325 3.2850 0.8925 ;
        RECT 3.1200 0.4875 3.1800 0.5475 ;
        RECT 3.0150 0.1275 3.0750 0.1875 ;
        RECT 3.0150 0.6825 3.0750 0.7425 ;
        RECT 2.9100 0.4875 2.9700 0.5475 ;
        RECT 2.8050 0.3075 2.8650 0.3675 ;
        RECT 2.8050 0.8325 2.8650 0.8925 ;
        RECT 2.7000 0.4875 2.7600 0.5475 ;
        RECT 2.5950 0.1425 2.6550 0.2025 ;
        RECT 2.5950 0.6825 2.6550 0.7425 ;
        RECT 2.4900 0.4875 2.5500 0.5475 ;
        RECT 2.3850 0.3075 2.4450 0.3675 ;
        RECT 2.3850 0.8325 2.4450 0.8925 ;
        RECT 2.2800 0.4875 2.3400 0.5475 ;
        RECT 2.1750 0.1425 2.2350 0.2025 ;
        RECT 2.1750 0.6825 2.2350 0.7425 ;
        RECT 2.0700 0.4875 2.1300 0.5475 ;
        RECT 1.9650 0.3075 2.0250 0.3675 ;
        RECT 1.9650 0.8325 2.0250 0.8925 ;
        RECT 1.8600 0.4875 1.9200 0.5475 ;
        RECT 1.7550 0.1425 1.8150 0.2025 ;
        RECT 1.7550 0.7575 1.8150 0.8175 ;
        RECT 1.6500 0.4875 1.7100 0.5475 ;
        RECT 1.5450 0.3075 1.6050 0.3675 ;
        RECT 1.5450 0.6675 1.6050 0.7275 ;
        RECT 1.4400 0.4875 1.5000 0.5475 ;
        RECT 1.3350 0.1425 1.3950 0.2025 ;
        RECT 1.3350 0.8325 1.3950 0.8925 ;
        RECT 1.2300 0.4875 1.2900 0.5475 ;
        RECT 1.1250 0.3075 1.1850 0.3675 ;
        RECT 1.1250 0.6675 1.1850 0.7275 ;
        RECT 1.0200 0.4875 1.0800 0.5475 ;
        RECT 0.9150 0.1425 0.9750 0.2025 ;
        RECT 0.9150 0.8325 0.9750 0.8925 ;
        RECT 0.8100 0.4875 0.8700 0.5475 ;
        RECT 0.7050 0.3075 0.7650 0.3675 ;
        RECT 0.7050 0.6675 0.7650 0.7275 ;
        RECT 0.6000 0.4875 0.6600 0.5475 ;
        RECT 0.4950 0.1425 0.5550 0.2025 ;
        RECT 0.4950 0.8325 0.5550 0.8925 ;
        RECT 0.3900 0.4875 0.4500 0.5475 ;
        RECT 0.2850 0.3075 0.3450 0.3675 ;
        RECT 0.2850 0.6675 0.3450 0.7275 ;
        RECT 0.1800 0.4875 0.2400 0.5475 ;
        RECT 0.0750 0.1575 0.1350 0.2175 ;
        RECT 0.0750 0.8175 0.1350 0.8775 ;
        LAYER M1 ;
        RECT 6.9975 0.6675 7.0725 0.8250 ;
        RECT 3.6900 0.6675 6.9975 0.7425 ;
        RECT 5.4000 0.4575 6.9675 0.5775 ;
        RECT 6.7725 0.2550 6.8775 0.3825 ;
        RECT 0.2550 0.3075 6.7725 0.3825 ;
        RECT 3.7425 0.4575 5.3100 0.5775 ;
        RECT 1.9275 0.8250 5.2425 0.9000 ;
        RECT 3.6150 0.6375 3.6900 0.7425 ;
        RECT 3.4350 0.6450 3.5325 0.7500 ;
        RECT 1.8225 0.6750 3.4350 0.7500 ;
        RECT 1.8525 0.4575 3.3975 0.5775 ;
        RECT 1.7475 0.6750 1.8225 0.9000 ;
        RECT 0.1575 0.8250 1.7475 0.9000 ;
        RECT 0.2625 0.6450 1.6350 0.7500 ;
        RECT 0.0525 0.7950 0.1575 0.9000 ;
    END
END NR4_0111


MACRO NR4_1000
    CLASS CORE ;
    FOREIGN NR4_1000 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.0500 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.9375 0.3075 1.0125 0.9000 ;
        RECT 0.7875 0.3075 0.9375 0.3825 ;
        RECT 0.9075 0.6675 0.9375 0.9000 ;
        RECT 0.6750 0.1500 0.7875 0.3825 ;
        RECT 0.3675 0.2550 0.6750 0.3375 ;
        RECT 0.2625 0.1500 0.3675 0.3375 ;
        END
    END ZN
    PIN A4
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1425 0.4500 0.2325 0.6000 ;
        RECT 0.0675 0.3675 0.1425 0.6825 ;
        END
    END A4
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.4125 0.4125 0.4725 0.5625 ;
        RECT 0.3075 0.4125 0.4125 0.7275 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.4125 0.8625 0.9600 0.9375 ;
        RECT 0.2475 0.8175 0.4125 0.9375 ;
        VIA 0.3300 0.8550 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.6975 0.5625 0.8925 0.6375 ;
        RECT 0.6225 0.1125 0.6975 0.6375 ;
        RECT 0.1050 0.1125 0.6225 0.1875 ;
        VIA 0.7950 0.6000 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.0050 -0.0750 1.0500 0.0750 ;
        RECT 0.8850 -0.0750 1.0050 0.2175 ;
        RECT 0.5850 -0.0750 0.8850 0.0750 ;
        RECT 0.4650 -0.0750 0.5850 0.1800 ;
        RECT 0.1425 -0.0750 0.4650 0.0750 ;
        RECT 0.0675 -0.0750 0.1425 0.2475 ;
        RECT 0.0000 -0.0750 0.0675 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.1425 0.9750 1.0500 1.1250 ;
        RECT 0.0675 0.8025 0.1425 1.1250 ;
        RECT 0.0000 0.9750 0.0675 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 0.9150 0.1575 0.9750 0.2175 ;
        RECT 0.9150 0.7575 0.9750 0.8175 ;
        RECT 0.8025 0.4950 0.8625 0.5550 ;
        RECT 0.7050 0.1725 0.7650 0.2325 ;
        RECT 0.5925 0.4950 0.6525 0.5550 ;
        RECT 0.4950 0.1200 0.5550 0.1800 ;
        RECT 0.3825 0.4800 0.4425 0.5400 ;
        RECT 0.2850 0.1725 0.3450 0.2325 ;
        RECT 0.1725 0.4950 0.2325 0.5550 ;
        RECT 0.0750 0.1575 0.1350 0.2175 ;
        RECT 0.0750 0.8325 0.1350 0.8925 ;
        LAYER M1 ;
        RECT 0.8325 0.4575 0.8625 0.5925 ;
        RECT 0.7575 0.4575 0.8325 0.8325 ;
        RECT 0.6225 0.4575 0.6525 0.5925 ;
        RECT 0.5475 0.4575 0.6225 0.9000 ;
        RECT 0.2475 0.8175 0.5475 0.9000 ;
    END
END NR4_1000


MACRO NR4_1010
    CLASS CORE ;
    FOREIGN NR4_1010 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.8900 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 0.7725 0.7125 1.2375 0.7875 ;
        RECT 0.7725 0.2625 0.8625 0.3375 ;
        RECT 0.6975 0.2625 0.7725 0.7875 ;
        VIA 0.9600 0.7500 VIA12_square ;
        VIA 0.7800 0.3000 VIA12_square ;
        END
    END ZN
    PIN A4
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.0725 0.4125 1.5375 0.4875 ;
        VIA 1.3650 0.4500 VIA12_square ;
        END
    END A4
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.7475 0.3675 1.8225 0.5325 ;
        RECT 1.7175 0.4200 1.7475 0.5325 ;
        RECT 1.6425 0.4200 1.7175 0.7200 ;
        RECT 1.1475 0.6450 1.6425 0.7200 ;
        RECT 1.0725 0.4350 1.1475 0.7200 ;
        RECT 1.0125 0.4350 1.0725 0.5550 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.8400 0.4350 0.8775 0.5550 ;
        RECT 0.7650 0.4350 0.8400 0.7200 ;
        RECT 0.2400 0.6450 0.7650 0.7200 ;
        RECT 0.1650 0.4350 0.2400 0.7200 ;
        RECT 0.1425 0.4350 0.1650 0.5325 ;
        RECT 0.0675 0.3675 0.1425 0.5325 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.5625 0.1125 1.0275 0.1875 ;
        RECT 0.4875 0.1125 0.5625 0.5850 ;
        VIA 0.5250 0.5025 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.8375 -0.0750 1.8900 0.0750 ;
        RECT 1.7325 -0.0750 1.8375 0.2400 ;
        RECT 1.4250 -0.0750 1.7325 0.0750 ;
        RECT 1.3050 -0.0750 1.4250 0.1875 ;
        RECT 1.0050 -0.0750 1.3050 0.0750 ;
        RECT 0.8850 -0.0750 1.0050 0.1875 ;
        RECT 0.5850 -0.0750 0.8850 0.0750 ;
        RECT 0.4650 -0.0750 0.5850 0.1875 ;
        RECT 0.1575 -0.0750 0.4650 0.0750 ;
        RECT 0.0525 -0.0750 0.1575 0.2400 ;
        RECT 0.0000 -0.0750 0.0525 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.4175 0.9750 1.8900 1.1250 ;
        RECT 1.3125 0.8325 1.4175 1.1250 ;
        RECT 0.0000 0.9750 1.3125 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.7550 0.1575 1.8150 0.2175 ;
        RECT 1.7550 0.8175 1.8150 0.8775 ;
        RECT 1.6500 0.4650 1.7100 0.5250 ;
        RECT 1.5450 0.1725 1.6050 0.2325 ;
        RECT 1.4400 0.4575 1.5000 0.5175 ;
        RECT 1.3350 0.1200 1.3950 0.1800 ;
        RECT 1.3350 0.8625 1.3950 0.9225 ;
        RECT 1.2300 0.4575 1.2900 0.5175 ;
        RECT 1.1250 0.1725 1.1850 0.2325 ;
        RECT 1.0200 0.4650 1.0800 0.5250 ;
        RECT 0.9150 0.1200 0.9750 0.1800 ;
        RECT 0.8100 0.4650 0.8700 0.5250 ;
        RECT 0.7050 0.1725 0.7650 0.2325 ;
        RECT 0.6000 0.4650 0.6600 0.5250 ;
        RECT 0.4950 0.1200 0.5550 0.1800 ;
        RECT 0.2850 0.1725 0.3450 0.2325 ;
        RECT 0.1800 0.4650 0.2400 0.5250 ;
        RECT 0.0750 0.1575 0.1350 0.2175 ;
        RECT 0.0750 0.8175 0.1350 0.8775 ;
        RECT 0.4950 0.8175 0.5550 0.8775 ;
        RECT 0.3900 0.4650 0.4500 0.5250 ;
        LAYER M1 ;
        RECT 1.4925 0.7950 1.8375 0.9000 ;
        RECT 1.5225 0.1500 1.6275 0.3375 ;
        RECT 1.2225 0.4125 1.5300 0.5550 ;
        RECT 1.2075 0.2625 1.5225 0.3375 ;
        RECT 1.1025 0.1500 1.2075 0.3375 ;
        RECT 0.7875 0.2625 1.1025 0.3375 ;
        RECT 0.9225 0.6675 0.9975 0.9000 ;
        RECT 0.4725 0.7950 0.9225 0.9000 ;
        RECT 0.6825 0.1500 0.7875 0.3375 ;
        RECT 0.3675 0.2625 0.6825 0.3375 ;
        RECT 0.3150 0.4200 0.6600 0.5700 ;
        RECT 0.2550 0.1500 0.3675 0.3375 ;
        RECT 0.0525 0.7950 0.3675 0.9000 ;
        LAYER VIA1 ;
        RECT 1.5375 0.8100 1.6125 0.8850 ;
        RECT 0.2475 0.8100 0.3225 0.8850 ;
        LAYER M2 ;
        RECT 1.5375 0.7650 1.6125 0.9375 ;
        RECT 0.3225 0.8625 1.5375 0.9375 ;
        RECT 0.2475 0.7650 0.3225 0.9375 ;
    END
END NR4_1010


MACRO OA211_0011
    CLASS CORE ;
    FOREIGN OA211_0011 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.4700 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 1.3575 0.3075 1.4325 0.7425 ;
        RECT 1.1925 0.3075 1.3575 0.3825 ;
        RECT 1.1925 0.6675 1.3575 0.7425 ;
        RECT 1.1175 0.2175 1.1925 0.3825 ;
        RECT 1.1175 0.6675 1.1925 0.8550 ;
        END
    END Z
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.8325 0.2625 1.1925 0.3375 ;
        RECT 0.7275 0.2325 0.8325 0.3375 ;
        VIA 0.9075 0.3000 VIA12_square ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.7575 0.8625 1.1925 0.9375 ;
        RECT 0.6525 0.4800 0.7575 0.9375 ;
        VIA 0.7050 0.5625 VIA12_square ;
        END
    END B
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1725 0.4575 0.2400 0.6000 ;
        RECT 0.1425 0.4575 0.1725 0.6975 ;
        RECT 0.0675 0.3675 0.1425 0.6975 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.4275 0.1125 0.6075 0.1875 ;
        RECT 0.3525 0.1125 0.4275 0.6450 ;
        RECT 0.0675 0.1125 0.3525 0.1875 ;
        VIA 0.3900 0.5325 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.4250 -0.0750 1.4700 0.0750 ;
        RECT 1.3050 -0.0750 1.4250 0.2175 ;
        RECT 1.0050 -0.0750 1.3050 0.0750 ;
        RECT 0.8850 -0.0750 1.0050 0.1875 ;
        RECT 0.0000 -0.0750 0.8850 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.4250 0.9750 1.4700 1.1250 ;
        RECT 1.3050 0.8175 1.4250 1.1250 ;
        RECT 1.0050 0.9750 1.3050 1.1250 ;
        RECT 0.8850 0.8700 1.0050 1.1250 ;
        RECT 0.5850 0.9750 0.8850 1.1250 ;
        RECT 0.4650 0.8700 0.5850 1.1250 ;
        RECT 0.0000 0.9750 0.4650 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.3350 0.1575 1.3950 0.2175 ;
        RECT 1.3350 0.8325 1.3950 0.8925 ;
        RECT 1.2225 0.4950 1.2825 0.5550 ;
        RECT 1.1250 0.2775 1.1850 0.3375 ;
        RECT 1.1250 0.7650 1.1850 0.8250 ;
        RECT 1.0200 0.4950 1.0800 0.5550 ;
        RECT 0.9150 0.1200 0.9750 0.1800 ;
        RECT 0.9150 0.8700 0.9750 0.9300 ;
        RECT 0.8175 0.4950 0.8775 0.5550 ;
        RECT 0.7050 0.7275 0.7650 0.7875 ;
        RECT 0.6000 0.4950 0.6600 0.5550 ;
        RECT 0.4950 0.1575 0.5550 0.2175 ;
        RECT 0.4950 0.8700 0.5550 0.9300 ;
        RECT 0.3900 0.4950 0.4500 0.5550 ;
        RECT 0.2850 0.3075 0.3450 0.3675 ;
        RECT 0.1800 0.4950 0.2400 0.5550 ;
        RECT 0.0750 0.1800 0.1350 0.2400 ;
        RECT 0.0750 0.8025 0.1350 0.8625 ;
        LAYER M1 ;
        RECT 1.0425 0.4650 1.2825 0.5850 ;
        RECT 0.9675 0.4650 1.0425 0.7950 ;
        RECT 0.8925 0.2625 0.9900 0.3675 ;
        RECT 0.3600 0.7200 0.9675 0.7950 ;
        RECT 0.8175 0.2625 0.8925 0.6150 ;
        RECT 0.5625 0.4500 0.7425 0.6450 ;
        RECT 0.2475 0.3000 0.6750 0.3750 ;
        RECT 0.1425 0.1500 0.5925 0.2250 ;
        RECT 0.3150 0.4500 0.4800 0.6450 ;
        RECT 0.2850 0.7200 0.3600 0.8850 ;
        RECT 0.0525 0.7800 0.2850 0.8850 ;
        RECT 0.0675 0.1500 0.1425 0.2700 ;
        LAYER VIA1 ;
        RECT 0.5325 0.3000 0.6075 0.3750 ;
        RECT 0.5025 0.7200 0.5775 0.7950 ;
        LAYER M2 ;
        RECT 0.5775 0.2700 0.6375 0.4050 ;
        RECT 0.5025 0.2700 0.5775 0.8400 ;
    END
END OA211_0011


MACRO OA211_0111
    CLASS CORE ;
    FOREIGN OA211_0111 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.9400 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 2.2575 0.2550 2.5725 0.7650 ;
        VIA 2.4150 0.3375 VIA12_slot ;
        VIA 2.4150 0.6825 VIA12_slot ;
        END
    END Z
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.7850 0.4350 1.8900 0.7875 ;
        RECT 1.3200 0.7125 1.7850 0.7875 ;
        RECT 1.2150 0.4350 1.3200 0.7875 ;
        VIA 1.8375 0.5325 VIA12_square ;
        VIA 1.2675 0.5175 VIA12_square ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.5300 0.2625 1.6350 0.5925 ;
        RECT 1.0800 0.2625 1.5300 0.3375 ;
        VIA 1.5825 0.5100 VIA12_square ;
        END
    END B
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.7725 0.4650 0.8775 0.7875 ;
        RECT 0.4425 0.7125 0.7725 0.7875 ;
        RECT 0.3675 0.5625 0.4425 0.7875 ;
        RECT 0.1500 0.5625 0.3675 0.6375 ;
        VIA 0.8250 0.5550 VIA12_square ;
        VIA 0.2325 0.6000 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.5175 0.2625 0.6225 0.5925 ;
        RECT 0.0900 0.2625 0.5175 0.3375 ;
        VIA 0.5700 0.5100 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 2.8875 -0.0750 2.9400 0.0750 ;
        RECT 2.7825 -0.0750 2.8875 0.3075 ;
        RECT 2.4750 -0.0750 2.7825 0.0750 ;
        RECT 2.3550 -0.0750 2.4750 0.1950 ;
        RECT 2.0550 -0.0750 2.3550 0.0750 ;
        RECT 1.9350 -0.0750 2.0550 0.1875 ;
        RECT 1.2150 -0.0750 1.9350 0.0750 ;
        RECT 1.0950 -0.0750 1.2150 0.2250 ;
        RECT 0.0000 -0.0750 1.0950 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 2.8875 0.9750 2.9400 1.1250 ;
        RECT 2.7825 0.6450 2.8875 1.1250 ;
        RECT 2.4750 0.9750 2.7825 1.1250 ;
        RECT 2.3550 0.8250 2.4750 1.1250 ;
        RECT 2.0550 0.9750 2.3550 1.1250 ;
        RECT 1.9350 0.8625 2.0550 1.1250 ;
        RECT 1.6350 0.9750 1.9350 1.1250 ;
        RECT 1.5150 0.8625 1.6350 1.1250 ;
        RECT 1.2075 0.9750 1.5150 1.1250 ;
        RECT 1.1025 0.8100 1.2075 1.1250 ;
        RECT 0.5850 0.9750 1.1025 1.1250 ;
        RECT 0.4650 0.8625 0.5850 1.1250 ;
        RECT 0.0000 0.9750 0.4650 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 2.8050 0.2175 2.8650 0.2775 ;
        RECT 2.8050 0.6675 2.8650 0.7275 ;
        RECT 2.8050 0.8325 2.8650 0.8925 ;
        RECT 2.7000 0.4800 2.7600 0.5400 ;
        RECT 2.5950 0.3075 2.6550 0.3675 ;
        RECT 2.5950 0.6525 2.6550 0.7125 ;
        RECT 2.4900 0.4800 2.5500 0.5400 ;
        RECT 2.3850 0.1275 2.4450 0.1875 ;
        RECT 2.3850 0.8325 2.4450 0.8925 ;
        RECT 2.2800 0.4800 2.3400 0.5400 ;
        RECT 2.1750 0.3075 2.2350 0.3675 ;
        RECT 2.1750 0.6525 2.2350 0.7125 ;
        RECT 2.0700 0.4800 2.1300 0.5400 ;
        RECT 1.9650 0.1275 2.0250 0.1875 ;
        RECT 1.9650 0.8625 2.0250 0.9225 ;
        RECT 1.8600 0.4950 1.9200 0.5550 ;
        RECT 1.7550 0.7200 1.8150 0.7800 ;
        RECT 1.6500 0.4800 1.7100 0.5400 ;
        RECT 1.5450 0.3000 1.6050 0.3600 ;
        RECT 1.5450 0.8625 1.6050 0.9225 ;
        RECT 1.4400 0.4800 1.5000 0.5400 ;
        RECT 1.3350 0.6600 1.3950 0.7200 ;
        RECT 1.2300 0.4800 1.2900 0.5400 ;
        RECT 1.1250 0.1575 1.1850 0.2175 ;
        RECT 1.1250 0.8325 1.1850 0.8925 ;
        RECT 0.9150 0.3075 0.9750 0.3675 ;
        RECT 0.9150 0.7200 0.9750 0.7800 ;
        RECT 0.8100 0.4950 0.8700 0.5550 ;
        RECT 0.7050 0.1650 0.7650 0.2250 ;
        RECT 0.6000 0.4800 0.6600 0.5400 ;
        RECT 0.4950 0.3075 0.5550 0.3675 ;
        RECT 0.4950 0.8625 0.5550 0.9225 ;
        RECT 0.3900 0.4800 0.4500 0.5400 ;
        RECT 0.2850 0.1650 0.3450 0.2250 ;
        RECT 0.1800 0.4800 0.2400 0.5400 ;
        RECT 0.0750 0.2925 0.1350 0.3525 ;
        RECT 0.0750 0.7425 0.1350 0.8025 ;
        LAYER M1 ;
        RECT 2.0775 0.4725 2.7900 0.5475 ;
        RECT 2.1525 0.2775 2.6850 0.3975 ;
        RECT 2.1525 0.6225 2.6850 0.7425 ;
        RECT 2.0025 0.4725 2.0775 0.7875 ;
        RECT 1.5300 0.7125 2.0025 0.7875 ;
        RECT 1.7850 0.3975 1.9275 0.6375 ;
        RECT 1.4325 0.4500 1.7100 0.5700 ;
        RECT 1.0500 0.3000 1.6650 0.3750 ;
        RECT 1.4550 0.6450 1.5300 0.7875 ;
        RECT 1.0275 0.6450 1.4550 0.7200 ;
        RECT 1.0950 0.4500 1.3575 0.5700 ;
        RECT 0.9975 0.3000 1.0500 0.3825 ;
        RECT 0.9525 0.6450 1.0275 0.7875 ;
        RECT 0.7575 0.3075 0.9975 0.3825 ;
        RECT 0.8775 0.4650 0.9900 0.5700 ;
        RECT 0.7950 0.1500 0.9600 0.2325 ;
        RECT 0.1575 0.7125 0.9525 0.7875 ;
        RECT 0.7350 0.4650 0.8775 0.6375 ;
        RECT 0.2550 0.1500 0.7950 0.2250 ;
        RECT 0.7200 0.3000 0.7575 0.3825 ;
        RECT 0.1575 0.3000 0.7200 0.3750 ;
        RECT 0.3900 0.4500 0.6600 0.5700 ;
        RECT 0.1200 0.4500 0.3150 0.6375 ;
        RECT 0.0525 0.2700 0.1575 0.3750 ;
        RECT 0.0525 0.7125 0.1575 0.8250 ;
        LAYER VIA1 ;
        RECT 2.0025 0.5175 2.0775 0.5925 ;
        RECT 0.8400 0.1575 0.9150 0.2325 ;
        LAYER M2 ;
        RECT 1.9875 0.1125 2.0925 0.6375 ;
        RECT 0.9600 0.1125 1.9875 0.1875 ;
        RECT 0.7950 0.1125 0.9600 0.2325 ;
    END
END OA211_0111


MACRO OA211_1000
    CLASS CORE ;
    FOREIGN OA211_1000 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.2600 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 1.1475 0.1500 1.2225 0.9000 ;
        RECT 1.1175 0.1500 1.1475 0.3825 ;
        RECT 1.1175 0.6675 1.1475 0.9000 ;
        END
    END Z
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.8325 0.2625 1.1925 0.3375 ;
        RECT 0.7275 0.2325 0.8325 0.3375 ;
        VIA 0.9075 0.3000 VIA12_square ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.7575 0.8625 1.1925 0.9375 ;
        RECT 0.6525 0.4800 0.7575 0.9375 ;
        VIA 0.7050 0.5625 VIA12_square ;
        END
    END B
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1725 0.4575 0.2400 0.6000 ;
        RECT 0.1425 0.4575 0.1725 0.6975 ;
        RECT 0.0675 0.3675 0.1425 0.6975 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.4275 0.1125 0.6075 0.1875 ;
        RECT 0.3525 0.1125 0.4275 0.6450 ;
        RECT 0.0675 0.1125 0.3525 0.1875 ;
        VIA 0.3900 0.5325 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.0050 -0.0750 1.2600 0.0750 ;
        RECT 0.8850 -0.0750 1.0050 0.1875 ;
        RECT 0.0000 -0.0750 0.8850 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.0050 0.9750 1.2600 1.1250 ;
        RECT 0.8850 0.8700 1.0050 1.1250 ;
        RECT 0.5850 0.9750 0.8850 1.1250 ;
        RECT 0.4650 0.8700 0.5850 1.1250 ;
        RECT 0.0000 0.9750 0.4650 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.1250 0.1800 1.1850 0.2400 ;
        RECT 1.1250 0.8100 1.1850 0.8700 ;
        RECT 1.0125 0.4950 1.0725 0.5550 ;
        RECT 0.9150 0.1200 0.9750 0.1800 ;
        RECT 0.9150 0.8700 0.9750 0.9300 ;
        RECT 0.8175 0.4950 0.8775 0.5550 ;
        RECT 0.7050 0.7950 0.7650 0.8550 ;
        RECT 0.6000 0.4950 0.6600 0.5550 ;
        RECT 0.4950 0.1575 0.5550 0.2175 ;
        RECT 0.4950 0.8700 0.5550 0.9300 ;
        RECT 0.3900 0.4950 0.4500 0.5550 ;
        RECT 0.2850 0.3075 0.3450 0.3675 ;
        RECT 0.1800 0.4950 0.2400 0.5550 ;
        RECT 0.0750 0.1800 0.1350 0.2400 ;
        RECT 0.0750 0.8100 0.1350 0.8700 ;
        LAYER M1 ;
        RECT 1.0425 0.4650 1.0725 0.5850 ;
        RECT 0.9675 0.4650 1.0425 0.7950 ;
        RECT 0.8925 0.2625 0.9900 0.3675 ;
        RECT 0.7875 0.7200 0.9675 0.7950 ;
        RECT 0.8175 0.2625 0.8925 0.6150 ;
        RECT 0.6825 0.7200 0.7875 0.8775 ;
        RECT 0.5625 0.4500 0.7425 0.6450 ;
        RECT 0.3600 0.7200 0.6825 0.7950 ;
        RECT 0.2475 0.3000 0.6750 0.3750 ;
        RECT 0.1425 0.1500 0.5925 0.2250 ;
        RECT 0.3150 0.4500 0.4800 0.6450 ;
        RECT 0.2850 0.7200 0.3600 0.8925 ;
        RECT 0.0525 0.7875 0.2850 0.8925 ;
        RECT 0.0675 0.1500 0.1425 0.2700 ;
        LAYER VIA1 ;
        RECT 0.5325 0.3000 0.6075 0.3750 ;
        RECT 0.5025 0.7200 0.5775 0.7950 ;
        LAYER M2 ;
        RECT 0.5775 0.2700 0.6375 0.4050 ;
        RECT 0.5025 0.2700 0.5775 0.8400 ;
    END
END OA211_1000


MACRO OA211_1010
    CLASS CORE ;
    FOREIGN OA211_1010 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.2600 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 1.1475 0.2175 1.2225 0.8325 ;
        RECT 1.1175 0.2175 1.1475 0.3825 ;
        RECT 1.1175 0.6675 1.1475 0.8325 ;
        END
    END Z
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.8325 0.2625 1.1925 0.3375 ;
        RECT 0.7275 0.2325 0.8325 0.3375 ;
        VIA 0.9075 0.3000 VIA12_square ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.7575 0.8625 1.1925 0.9375 ;
        RECT 0.6525 0.4800 0.7575 0.9375 ;
        VIA 0.7050 0.5625 VIA12_square ;
        END
    END B
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1725 0.4575 0.2400 0.6000 ;
        RECT 0.1425 0.4575 0.1725 0.6975 ;
        RECT 0.0675 0.3675 0.1425 0.6975 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.4275 0.1125 0.6075 0.1875 ;
        RECT 0.3525 0.1125 0.4275 0.6450 ;
        RECT 0.0675 0.1125 0.3525 0.1875 ;
        VIA 0.3900 0.5325 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.0050 -0.0750 1.2600 0.0750 ;
        RECT 0.8850 -0.0750 1.0050 0.1875 ;
        RECT 0.0000 -0.0750 0.8850 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.0050 0.9750 1.2600 1.1250 ;
        RECT 0.8850 0.8700 1.0050 1.1250 ;
        RECT 0.5850 0.9750 0.8850 1.1250 ;
        RECT 0.4650 0.8700 0.5850 1.1250 ;
        RECT 0.0000 0.9750 0.4650 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.1250 0.2700 1.1850 0.3300 ;
        RECT 1.1250 0.7200 1.1850 0.7800 ;
        RECT 1.0125 0.4950 1.0725 0.5550 ;
        RECT 0.9150 0.1200 0.9750 0.1800 ;
        RECT 0.9150 0.8700 0.9750 0.9300 ;
        RECT 0.8175 0.4950 0.8775 0.5550 ;
        RECT 0.7050 0.7275 0.7650 0.7875 ;
        RECT 0.6000 0.4950 0.6600 0.5550 ;
        RECT 0.4950 0.1575 0.5550 0.2175 ;
        RECT 0.4950 0.8700 0.5550 0.9300 ;
        RECT 0.3900 0.4950 0.4500 0.5550 ;
        RECT 0.2850 0.3075 0.3450 0.3675 ;
        RECT 0.1800 0.4950 0.2400 0.5550 ;
        RECT 0.0750 0.1800 0.1350 0.2400 ;
        RECT 0.0750 0.8025 0.1350 0.8625 ;
        LAYER M1 ;
        RECT 1.0425 0.4650 1.0725 0.5850 ;
        RECT 0.9675 0.4650 1.0425 0.7950 ;
        RECT 0.8925 0.2625 0.9900 0.3675 ;
        RECT 0.3600 0.7200 0.9675 0.7950 ;
        RECT 0.8175 0.2625 0.8925 0.6150 ;
        RECT 0.5625 0.4500 0.7425 0.6450 ;
        RECT 0.2475 0.3000 0.6750 0.3750 ;
        RECT 0.1425 0.1500 0.5925 0.2250 ;
        RECT 0.3150 0.4500 0.4800 0.6450 ;
        RECT 0.2850 0.7200 0.3600 0.8850 ;
        RECT 0.0525 0.7800 0.2850 0.8850 ;
        RECT 0.0675 0.1500 0.1425 0.2700 ;
        LAYER VIA1 ;
        RECT 0.5325 0.3000 0.6075 0.3750 ;
        RECT 0.5025 0.7200 0.5775 0.7950 ;
        LAYER M2 ;
        RECT 0.5775 0.2700 0.6375 0.4050 ;
        RECT 0.5025 0.2700 0.5775 0.8400 ;
    END
END OA211_1010


MACRO OA21_0011
    CLASS CORE ;
    FOREIGN OA21_0011 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.2600 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 1.1475 0.3075 1.2225 0.7425 ;
        RECT 0.9825 0.3075 1.1475 0.3825 ;
        RECT 0.9825 0.6675 1.1475 0.7425 ;
        RECT 0.9075 0.2175 0.9825 0.3825 ;
        RECT 0.9075 0.6675 0.9825 0.8550 ;
        END
    END Z
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.5175 0.5625 0.9825 0.6375 ;
        VIA 0.6000 0.6000 VIA12_square ;
        END
    END B
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1425 0.4650 0.2325 0.6825 ;
        RECT 0.0675 0.3675 0.1425 0.6825 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.2025 0.7125 0.6675 0.7875 ;
        VIA 0.3525 0.7500 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.2150 -0.0750 1.2600 0.0750 ;
        RECT 1.0950 -0.0750 1.2150 0.2175 ;
        RECT 0.7950 -0.0750 1.0950 0.0750 ;
        RECT 0.6900 -0.0750 0.7950 0.2250 ;
        RECT 0.0000 -0.0750 0.6900 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.2150 0.9750 1.2600 1.1250 ;
        RECT 1.0950 0.8175 1.2150 1.1250 ;
        RECT 0.7950 0.9750 1.0950 1.1250 ;
        RECT 0.6750 0.8700 0.7950 1.1250 ;
        RECT 0.1575 0.9750 0.6750 1.1250 ;
        RECT 0.0675 0.7950 0.1575 1.1250 ;
        RECT 0.0000 0.9750 0.0675 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.1250 0.1575 1.1850 0.2175 ;
        RECT 1.1250 0.8325 1.1850 0.8925 ;
        RECT 1.0125 0.4950 1.0725 0.5550 ;
        RECT 0.9150 0.2550 0.9750 0.3150 ;
        RECT 0.9150 0.7650 0.9750 0.8250 ;
        RECT 0.8025 0.4950 0.8625 0.5550 ;
        RECT 0.7050 0.1350 0.7650 0.1950 ;
        RECT 0.7050 0.8700 0.7650 0.9300 ;
        RECT 0.6000 0.4950 0.6600 0.5550 ;
        RECT 0.4950 0.1575 0.5550 0.2175 ;
        RECT 0.4950 0.7500 0.5550 0.8100 ;
        RECT 0.3825 0.4950 0.4425 0.5550 ;
        RECT 0.2850 0.3075 0.3450 0.3675 ;
        RECT 0.1725 0.4950 0.2325 0.5550 ;
        RECT 0.0750 0.1575 0.1350 0.2175 ;
        RECT 0.0750 0.8325 0.1350 0.8925 ;
        LAYER M1 ;
        RECT 0.8325 0.4650 1.0725 0.5850 ;
        RECT 0.7575 0.3000 0.8325 0.7950 ;
        RECT 0.2550 0.3000 0.7575 0.3750 ;
        RECT 0.5625 0.7200 0.7575 0.7950 ;
        RECT 0.5175 0.4500 0.6825 0.6450 ;
        RECT 0.4875 0.7200 0.5625 0.8400 ;
        RECT 0.3900 0.4650 0.4425 0.6300 ;
        RECT 0.3075 0.4650 0.3900 0.8325 ;
        RECT 0.0450 0.1500 0.1500 0.2550 ;
        RECT 0.1500 0.1500 0.5850 0.2250 ;
    END
END OA21_0011


MACRO OA21_0111
    CLASS CORE ;
    FOREIGN OA21_0111 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.3100 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 1.4175 0.2775 1.7325 0.7425 ;
        VIA 1.5750 0.3375 VIA12_slot ;
        VIA 1.5750 0.6825 VIA12_slot ;
        END
    END Z
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.9575 0.5625 2.2125 0.6375 ;
        RECT 1.8825 0.5625 1.9575 0.9375 ;
        RECT 1.0500 0.8625 1.8825 0.9375 ;
        RECT 0.9450 0.4425 1.0500 0.9375 ;
        VIA 2.1300 0.6000 VIA12_square ;
        VIA 0.9975 0.5250 VIA12_square ;
        END
    END B
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.5325 0.1125 0.6075 0.5850 ;
        RECT 0.0675 0.1125 0.5325 0.1875 ;
        VIA 0.5700 0.5025 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.8625 0.4650 0.8700 0.5850 ;
        RECT 0.7650 0.4650 0.8625 0.7050 ;
        RECT 0.2400 0.6300 0.7650 0.7050 ;
        RECT 0.1425 0.4650 0.2400 0.7050 ;
        RECT 0.0675 0.3675 0.1425 0.7050 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 2.0550 -0.0750 2.3100 0.0750 ;
        RECT 1.9350 -0.0750 2.0550 0.1800 ;
        RECT 1.6350 -0.0750 1.9350 0.0750 ;
        RECT 1.5150 -0.0750 1.6350 0.1950 ;
        RECT 1.1925 -0.0750 1.5150 0.0750 ;
        RECT 1.1175 -0.0750 1.1925 0.2100 ;
        RECT 0.0000 -0.0750 1.1175 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 2.0550 0.9750 2.3100 1.1250 ;
        RECT 1.9350 0.8700 2.0550 1.1250 ;
        RECT 1.6350 0.9750 1.9350 1.1250 ;
        RECT 1.5150 0.8625 1.6350 1.1250 ;
        RECT 1.2150 0.9750 1.5150 1.1250 ;
        RECT 1.0950 0.8700 1.2150 1.1250 ;
        RECT 0.5850 0.9750 1.0950 1.1250 ;
        RECT 0.4650 0.7800 0.5850 1.1250 ;
        RECT 0.0000 0.9750 0.4650 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 2.1750 0.2250 2.2350 0.2850 ;
        RECT 2.1750 0.7500 2.2350 0.8100 ;
        RECT 2.0700 0.4950 2.1300 0.5550 ;
        RECT 1.9650 0.1200 2.0250 0.1800 ;
        RECT 1.9650 0.8700 2.0250 0.9300 ;
        RECT 1.8600 0.4650 1.9200 0.5250 ;
        RECT 1.7550 0.2250 1.8150 0.2850 ;
        RECT 1.7550 0.7575 1.8150 0.8175 ;
        RECT 1.6500 0.4650 1.7100 0.5250 ;
        RECT 1.5450 0.1275 1.6050 0.1875 ;
        RECT 1.5450 0.8700 1.6050 0.9300 ;
        RECT 1.4400 0.4650 1.5000 0.5250 ;
        RECT 1.3350 0.2250 1.3950 0.2850 ;
        RECT 1.3350 0.7575 1.3950 0.8175 ;
        RECT 1.2300 0.4650 1.2900 0.5250 ;
        RECT 1.1250 0.1200 1.1850 0.1800 ;
        RECT 1.1250 0.8700 1.1850 0.9300 ;
        RECT 1.0200 0.4950 1.0800 0.5550 ;
        RECT 0.9150 0.1575 0.9750 0.2175 ;
        RECT 0.9150 0.8250 0.9750 0.8850 ;
        RECT 0.8100 0.4950 0.8700 0.5550 ;
        RECT 0.7050 0.3075 0.7650 0.3675 ;
        RECT 0.6000 0.4875 0.6600 0.5475 ;
        RECT 0.4950 0.1575 0.5550 0.2175 ;
        RECT 0.4950 0.8025 0.5550 0.8625 ;
        RECT 0.3900 0.4875 0.4500 0.5475 ;
        RECT 0.2850 0.3075 0.3450 0.3675 ;
        RECT 0.1800 0.4950 0.2400 0.5550 ;
        RECT 0.0750 0.1725 0.1350 0.2325 ;
        RECT 0.0750 0.8175 0.1350 0.8775 ;
        LAYER M1 ;
        RECT 2.1675 0.1875 2.2425 0.3600 ;
        RECT 2.0475 0.4350 2.2425 0.6450 ;
        RECT 2.1675 0.7200 2.2425 0.8400 ;
        RECT 1.8975 0.2550 2.1675 0.3600 ;
        RECT 1.9725 0.7200 2.1675 0.7950 ;
        RECT 1.8975 0.4575 1.9725 0.7950 ;
        RECT 1.2300 0.4575 1.8975 0.5475 ;
        RECT 1.7475 0.1950 1.8225 0.3825 ;
        RECT 1.7475 0.6225 1.8225 0.8700 ;
        RECT 1.4175 0.2925 1.7475 0.3825 ;
        RECT 1.4025 0.6225 1.7475 0.7425 ;
        RECT 1.3125 0.1950 1.4175 0.3825 ;
        RECT 1.3275 0.6225 1.4025 0.8700 ;
        RECT 1.1550 0.4575 1.2300 0.7950 ;
        RECT 1.0200 0.7200 1.1550 0.7950 ;
        RECT 0.9450 0.3900 1.0800 0.6450 ;
        RECT 0.9300 0.1500 1.0425 0.3150 ;
        RECT 0.9450 0.7200 1.0200 0.9000 ;
        RECT 0.6825 0.7950 0.9450 0.9000 ;
        RECT 0.1575 0.1500 0.9300 0.2250 ;
        RECT 0.2475 0.3000 0.8175 0.3750 ;
        RECT 0.3600 0.4500 0.6900 0.5550 ;
        RECT 0.0525 0.7950 0.3675 0.9000 ;
        RECT 0.0525 0.1500 0.1575 0.2550 ;
        LAYER VIA1 ;
        RECT 1.9425 0.2625 2.0175 0.3375 ;
        RECT 0.9375 0.1950 1.0125 0.2700 ;
        RECT 0.7275 0.7950 0.8025 0.8700 ;
        RECT 0.6975 0.3000 0.7725 0.3750 ;
        RECT 0.2475 0.7950 0.3225 0.8700 ;
        LAYER M2 ;
        RECT 1.9425 0.2625 2.0625 0.3375 ;
        RECT 1.8600 0.1125 1.9425 0.3375 ;
        RECT 1.0275 0.1125 1.8600 0.1875 ;
        RECT 0.9225 0.1125 1.0275 0.3150 ;
        RECT 0.7875 0.7800 0.8475 0.8850 ;
        RECT 0.6825 0.2625 0.7875 0.8850 ;
        RECT 0.1800 0.7950 0.6825 0.8850 ;
    END
END OA21_0111


MACRO OA21_1000
    CLASS CORE ;
    FOREIGN OA21_1000 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.0500 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.9375 0.1500 1.0125 0.9000 ;
        RECT 0.9075 0.1500 0.9375 0.3825 ;
        RECT 0.9075 0.6675 0.9375 0.9000 ;
        END
    END Z
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.5175 0.5625 0.9825 0.6375 ;
        VIA 0.6000 0.6000 VIA12_square ;
        END
    END B
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1425 0.4650 0.2325 0.6825 ;
        RECT 0.0675 0.3675 0.1425 0.6825 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.2025 0.7125 0.6675 0.7875 ;
        VIA 0.3525 0.7500 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.7950 -0.0750 1.0500 0.0750 ;
        RECT 0.6900 -0.0750 0.7950 0.2250 ;
        RECT 0.0000 -0.0750 0.6900 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.7950 0.9750 1.0500 1.1250 ;
        RECT 0.6750 0.8700 0.7950 1.1250 ;
        RECT 0.1575 0.9750 0.6750 1.1250 ;
        RECT 0.0675 0.7950 0.1575 1.1250 ;
        RECT 0.0000 0.9750 0.0675 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 0.9150 0.1800 0.9750 0.2400 ;
        RECT 0.9150 0.8100 0.9750 0.8700 ;
        RECT 0.8025 0.4950 0.8625 0.5550 ;
        RECT 0.7050 0.1350 0.7650 0.1950 ;
        RECT 0.7050 0.8700 0.7650 0.9300 ;
        RECT 0.6000 0.4950 0.6600 0.5550 ;
        RECT 0.4950 0.1575 0.5550 0.2175 ;
        RECT 0.4950 0.8025 0.5550 0.8625 ;
        RECT 0.3825 0.4950 0.4425 0.5550 ;
        RECT 0.2850 0.3075 0.3450 0.3675 ;
        RECT 0.1725 0.4950 0.2325 0.5550 ;
        RECT 0.0750 0.1575 0.1350 0.2175 ;
        RECT 0.0750 0.8325 0.1350 0.8925 ;
        LAYER M1 ;
        RECT 0.8325 0.4650 0.8625 0.5850 ;
        RECT 0.7575 0.3000 0.8325 0.7950 ;
        RECT 0.2550 0.3000 0.7575 0.3750 ;
        RECT 0.5775 0.7200 0.7575 0.7950 ;
        RECT 0.5175 0.4500 0.6825 0.6450 ;
        RECT 0.1500 0.1500 0.5850 0.2250 ;
        RECT 0.4725 0.7200 0.5775 0.8925 ;
        RECT 0.3900 0.4650 0.4425 0.6300 ;
        RECT 0.3075 0.4650 0.3900 0.8325 ;
        RECT 0.0450 0.1500 0.1500 0.2550 ;
    END
END OA21_1000


MACRO OA21_1010
    CLASS CORE ;
    FOREIGN OA21_1010 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.0500 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.9375 0.2175 1.0125 0.8325 ;
        RECT 0.9075 0.2175 0.9375 0.3825 ;
        RECT 0.9075 0.6675 0.9375 0.8325 ;
        END
    END Z
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.5175 0.5625 0.9825 0.6375 ;
        VIA 0.6000 0.6000 VIA12_square ;
        END
    END B
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1425 0.4650 0.2325 0.6825 ;
        RECT 0.0675 0.3675 0.1425 0.6825 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.2025 0.7125 0.6675 0.7875 ;
        VIA 0.3525 0.7500 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.7950 -0.0750 1.0500 0.0750 ;
        RECT 0.6900 -0.0750 0.7950 0.2250 ;
        RECT 0.0000 -0.0750 0.6900 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.7950 0.9750 1.0500 1.1250 ;
        RECT 0.6750 0.8700 0.7950 1.1250 ;
        RECT 0.1575 0.9750 0.6750 1.1250 ;
        RECT 0.0675 0.7950 0.1575 1.1250 ;
        RECT 0.0000 0.9750 0.0675 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 0.9150 0.2700 0.9750 0.3300 ;
        RECT 0.9150 0.7200 0.9750 0.7800 ;
        RECT 0.8025 0.4950 0.8625 0.5550 ;
        RECT 0.7050 0.1350 0.7650 0.1950 ;
        RECT 0.7050 0.8700 0.7650 0.9300 ;
        RECT 0.6000 0.4950 0.6600 0.5550 ;
        RECT 0.4950 0.1575 0.5550 0.2175 ;
        RECT 0.4950 0.7500 0.5550 0.8100 ;
        RECT 0.3825 0.4950 0.4425 0.5550 ;
        RECT 0.2850 0.3075 0.3450 0.3675 ;
        RECT 0.1725 0.4950 0.2325 0.5550 ;
        RECT 0.0750 0.1575 0.1350 0.2175 ;
        RECT 0.0750 0.8325 0.1350 0.8925 ;
        LAYER M1 ;
        RECT 0.8325 0.4650 0.8625 0.5850 ;
        RECT 0.7575 0.3000 0.8325 0.7950 ;
        RECT 0.2550 0.3000 0.7575 0.3750 ;
        RECT 0.5625 0.7200 0.7575 0.7950 ;
        RECT 0.5175 0.4500 0.6825 0.6450 ;
        RECT 0.1500 0.1500 0.5850 0.2250 ;
        RECT 0.4875 0.7200 0.5625 0.8400 ;
        RECT 0.3900 0.4650 0.4425 0.6300 ;
        RECT 0.3075 0.4650 0.3900 0.8325 ;
        RECT 0.0450 0.1500 0.1500 0.2550 ;
    END
END OA21_1010


MACRO OA221_0011
    CLASS CORE ;
    FOREIGN OA221_0011 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.8900 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 1.7775 0.3075 1.8525 0.7425 ;
        RECT 1.6125 0.3075 1.7775 0.3825 ;
        RECT 1.6125 0.6675 1.7775 0.7425 ;
        RECT 1.5375 0.2175 1.6125 0.3825 ;
        RECT 1.5375 0.6675 1.6125 0.8550 ;
        END
    END Z
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.1475 0.8625 1.6125 0.9375 ;
        RECT 1.0725 0.6000 1.1475 0.9375 ;
        RECT 0.7275 0.6000 1.0725 0.6750 ;
        RECT 0.6525 0.4875 0.7275 0.6750 ;
        VIA 0.6900 0.5700 VIA12_square ;
        END
    END C
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.1475 0.2625 1.6125 0.3375 ;
        RECT 1.1475 0.4125 1.2975 0.4875 ;
        RECT 1.0725 0.2625 1.1475 0.4875 ;
        VIA 1.2000 0.4500 VIA12_square ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.8775 0.1125 1.4175 0.1875 ;
        RECT 0.8775 0.4200 0.9675 0.5250 ;
        RECT 0.8025 0.1125 0.8775 0.5250 ;
        VIA 0.8850 0.4725 VIA12_square ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1425 0.4650 0.2475 0.5850 ;
        RECT 0.0675 0.3675 0.1425 0.6825 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.4275 0.1125 0.6075 0.1875 ;
        RECT 0.3525 0.1125 0.4275 0.6600 ;
        RECT 0.0675 0.1125 0.3525 0.1875 ;
        VIA 0.3900 0.5775 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.8450 -0.0750 1.8900 0.0750 ;
        RECT 1.7250 -0.0750 1.8450 0.2175 ;
        RECT 1.4250 -0.0750 1.7250 0.0750 ;
        RECT 1.3050 -0.0750 1.4250 0.3300 ;
        RECT 1.0050 -0.0750 1.3050 0.0750 ;
        RECT 0.8850 -0.0750 1.0050 0.1800 ;
        RECT 0.0000 -0.0750 0.8850 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.8450 0.9750 1.8900 1.1250 ;
        RECT 1.7250 0.8175 1.8450 1.1250 ;
        RECT 1.4250 0.9750 1.7250 1.1250 ;
        RECT 1.3050 0.8325 1.4250 1.1250 ;
        RECT 0.7650 0.9750 1.3050 1.1250 ;
        RECT 0.6600 0.8100 0.7650 1.1250 ;
        RECT 0.1650 0.9750 0.6600 1.1250 ;
        RECT 0.0450 0.8175 0.1650 1.1250 ;
        RECT 0.0000 0.9750 0.0450 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.7550 0.1575 1.8150 0.2175 ;
        RECT 1.7550 0.8325 1.8150 0.8925 ;
        RECT 1.6425 0.4950 1.7025 0.5550 ;
        RECT 1.5450 0.2775 1.6050 0.3375 ;
        RECT 1.5450 0.7650 1.6050 0.8250 ;
        RECT 1.4400 0.4950 1.5000 0.5550 ;
        RECT 1.3350 0.2400 1.3950 0.3000 ;
        RECT 1.3350 0.8325 1.3950 0.8925 ;
        RECT 1.1250 0.2325 1.1850 0.2925 ;
        RECT 1.1250 0.7725 1.1850 0.8325 ;
        RECT 1.0275 0.4950 1.0875 0.5550 ;
        RECT 0.9150 0.1200 0.9750 0.1800 ;
        RECT 0.8100 0.4950 0.8700 0.5550 ;
        RECT 0.7050 0.2325 0.7650 0.2925 ;
        RECT 0.7050 0.8400 0.7650 0.9000 ;
        RECT 0.6000 0.4950 0.6600 0.5550 ;
        RECT 0.4950 0.1575 0.5550 0.2175 ;
        RECT 0.4950 0.8100 0.5550 0.8700 ;
        RECT 0.3900 0.4950 0.4500 0.5550 ;
        RECT 0.2850 0.3150 0.3450 0.3750 ;
        RECT 0.1800 0.4950 0.2400 0.5550 ;
        RECT 0.0750 0.1650 0.1350 0.2250 ;
        RECT 0.0750 0.8325 0.1350 0.8925 ;
        LAYER M1 ;
        RECT 1.4625 0.4650 1.7025 0.5850 ;
        RECT 1.3875 0.4650 1.4625 0.7575 ;
        RECT 1.1925 0.6825 1.3875 0.7575 ;
        RECT 1.0275 0.4125 1.2975 0.6000 ;
        RECT 1.1175 0.6825 1.1925 0.8925 ;
        RECT 1.0950 0.1950 1.1850 0.3300 ;
        RECT 0.8400 0.7875 1.1175 0.8925 ;
        RECT 0.7950 0.2550 1.0950 0.3300 ;
        RECT 0.8100 0.4050 0.9525 0.6975 ;
        RECT 0.6975 0.2025 0.7950 0.3300 ;
        RECT 0.5700 0.4875 0.7275 0.7050 ;
        RECT 0.3825 0.3000 0.6225 0.4125 ;
        RECT 0.1500 0.1500 0.5850 0.2250 ;
        RECT 0.2775 0.7800 0.5850 0.8925 ;
        RECT 0.3300 0.4950 0.4950 0.7050 ;
        RECT 0.2550 0.3000 0.3825 0.3900 ;
        RECT 0.0450 0.1500 0.1500 0.2550 ;
        LAYER VIA1 ;
        RECT 0.8850 0.7875 0.9600 0.8625 ;
        RECT 0.5025 0.3375 0.5775 0.4125 ;
        RECT 0.4275 0.8175 0.5025 0.8925 ;
        LAYER M2 ;
        RECT 0.8400 0.7500 0.9900 0.8925 ;
        RECT 0.5775 0.7500 0.8400 0.8250 ;
        RECT 0.5775 0.2625 0.6075 0.3375 ;
        RECT 0.5025 0.2625 0.5775 0.8925 ;
        RECT 0.3825 0.8175 0.5025 0.8925 ;
    END
END OA221_0011


MACRO OA221_0111
    CLASS CORE ;
    FOREIGN OA221_0111 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.3600 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 2.6775 0.2400 2.9925 0.7500 ;
        VIA 2.8350 0.3225 VIA12_slot ;
        VIA 2.8350 0.6675 VIA12_slot ;
        END
    END Z
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.1025 0.1125 1.2075 0.6825 ;
        RECT 0.6375 0.1125 1.1025 0.1875 ;
        VIA 1.1550 0.5250 VIA12_square ;
        END
    END C
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 2.0475 0.2625 2.5200 0.3375 ;
        RECT 1.9425 0.2625 2.0475 0.6225 ;
        VIA 1.9950 0.5250 VIA12_square ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.6275 0.1125 2.0925 0.1875 ;
        RECT 1.5225 0.1125 1.6275 0.6900 ;
        VIA 1.5750 0.5775 VIA12_square ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.7725 0.4650 0.8775 0.7050 ;
        RECT 0.2400 0.6300 0.7725 0.7050 ;
        RECT 0.1425 0.4650 0.2400 0.7050 ;
        RECT 0.0675 0.3675 0.1425 0.7050 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.4725 0.4200 0.5775 0.7875 ;
        RECT 0.0900 0.7125 0.4725 0.7875 ;
        VIA 0.5250 0.5025 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 3.2925 -0.0750 3.3600 0.0750 ;
        RECT 3.2175 -0.0750 3.2925 0.3150 ;
        RECT 2.8950 -0.0750 3.2175 0.0750 ;
        RECT 2.7750 -0.0750 2.8950 0.1950 ;
        RECT 2.4525 -0.0750 2.7750 0.0750 ;
        RECT 2.3775 -0.0750 2.4525 0.3150 ;
        RECT 2.0550 -0.0750 2.3775 0.0750 ;
        RECT 1.9350 -0.0750 2.0550 0.2400 ;
        RECT 1.6350 -0.0750 1.9350 0.0750 ;
        RECT 1.5300 -0.0750 1.6350 0.2475 ;
        RECT 0.0000 -0.0750 1.5300 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 3.2925 0.9750 3.3600 1.1250 ;
        RECT 3.2175 0.6375 3.2925 1.1250 ;
        RECT 2.8725 0.9750 3.2175 1.1250 ;
        RECT 2.7975 0.8175 2.8725 1.1250 ;
        RECT 2.4750 0.9750 2.7975 1.1250 ;
        RECT 2.3550 0.8025 2.4750 1.1250 ;
        RECT 1.6350 0.9750 2.3550 1.1250 ;
        RECT 1.5150 0.8025 1.6350 1.1250 ;
        RECT 1.4175 0.9750 1.5150 1.1250 ;
        RECT 1.3125 0.6450 1.4175 1.1250 ;
        RECT 1.0125 0.9750 1.3125 1.1250 ;
        RECT 0.9150 0.8025 1.0125 1.1250 ;
        RECT 0.1575 0.9750 0.9150 1.1250 ;
        RECT 0.0525 0.8025 0.1575 1.1250 ;
        RECT 0.0000 0.9750 0.0525 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 3.2250 0.2250 3.2850 0.2850 ;
        RECT 3.2250 0.6675 3.2850 0.7275 ;
        RECT 3.2250 0.8325 3.2850 0.8925 ;
        RECT 3.1200 0.4650 3.1800 0.5250 ;
        RECT 3.0150 0.2250 3.0750 0.2850 ;
        RECT 3.0150 0.7575 3.0750 0.8175 ;
        RECT 2.9100 0.4650 2.9700 0.5250 ;
        RECT 2.8050 0.1275 2.8650 0.1875 ;
        RECT 2.8050 0.8475 2.8650 0.9075 ;
        RECT 2.7000 0.4650 2.7600 0.5250 ;
        RECT 2.5950 0.2250 2.6550 0.2850 ;
        RECT 2.5950 0.7575 2.6550 0.8175 ;
        RECT 2.4900 0.4650 2.5500 0.5250 ;
        RECT 2.3850 0.2100 2.4450 0.2700 ;
        RECT 2.3850 0.8250 2.4450 0.8850 ;
        RECT 2.2800 0.4950 2.3400 0.5550 ;
        RECT 2.1750 0.3225 2.2350 0.3825 ;
        RECT 2.0700 0.4950 2.1300 0.5550 ;
        RECT 1.9650 0.1500 2.0250 0.2100 ;
        RECT 1.9650 0.8175 2.0250 0.8775 ;
        RECT 1.8600 0.4950 1.9200 0.5550 ;
        RECT 1.7550 0.3225 1.8150 0.3825 ;
        RECT 1.6500 0.4950 1.7100 0.5550 ;
        RECT 1.5450 0.1575 1.6050 0.2175 ;
        RECT 1.5450 0.8175 1.6050 0.8775 ;
        RECT 1.3350 0.1575 1.3950 0.2175 ;
        RECT 1.3350 0.6675 1.3950 0.7275 ;
        RECT 1.3350 0.8325 1.3950 0.8925 ;
        RECT 1.2300 0.4950 1.2900 0.5550 ;
        RECT 1.1250 0.3225 1.1850 0.3825 ;
        RECT 1.1250 0.8100 1.1850 0.8700 ;
        RECT 1.0200 0.4950 1.0800 0.5550 ;
        RECT 0.9150 0.1575 0.9750 0.2175 ;
        RECT 0.9150 0.8325 0.9750 0.8925 ;
        RECT 0.8100 0.4950 0.8700 0.5550 ;
        RECT 0.7050 0.3075 0.7650 0.3675 ;
        RECT 0.6000 0.4800 0.6600 0.5400 ;
        RECT 0.4950 0.1575 0.5550 0.2175 ;
        RECT 0.4950 0.8025 0.5550 0.8625 ;
        RECT 0.3900 0.4800 0.4500 0.5400 ;
        RECT 0.2850 0.3075 0.3450 0.3675 ;
        RECT 0.1800 0.4950 0.2400 0.5550 ;
        RECT 0.0750 0.1725 0.1350 0.2325 ;
        RECT 0.0750 0.8325 0.1350 0.8925 ;
        LAYER M1 ;
        RECT 2.4900 0.4425 3.2100 0.5475 ;
        RECT 2.9925 0.1950 3.0975 0.3675 ;
        RECT 3.0075 0.6225 3.0825 0.8700 ;
        RECT 2.6625 0.6225 3.0075 0.7125 ;
        RECT 2.6775 0.2775 2.9925 0.3675 ;
        RECT 2.5725 0.1950 2.6775 0.3675 ;
        RECT 2.5875 0.6225 2.6625 0.8700 ;
        RECT 2.4150 0.4425 2.4900 0.6750 ;
        RECT 2.2350 0.4650 2.3400 0.7275 ;
        RECT 1.8525 0.3150 2.2650 0.3900 ;
        RECT 1.7325 0.6525 2.2350 0.7275 ;
        RECT 1.8225 0.8025 2.1675 0.9000 ;
        RECT 1.8300 0.4725 2.1525 0.5775 ;
        RECT 1.7175 0.3150 1.8525 0.3975 ;
        RECT 1.6575 0.4725 1.7325 0.7275 ;
        RECT 1.0950 0.3225 1.7175 0.3975 ;
        RECT 1.5375 0.4725 1.6575 0.6600 ;
        RECT 0.1575 0.1500 1.4250 0.2250 ;
        RECT 0.9900 0.4725 1.3200 0.5700 ;
        RECT 1.0875 0.6525 1.2375 0.8850 ;
        RECT 0.2475 0.3000 0.8925 0.3750 ;
        RECT 0.4650 0.7800 0.8400 0.8850 ;
        RECT 0.3600 0.4500 0.6900 0.5550 ;
        RECT 0.0525 0.1500 0.1575 0.2550 ;
        LAYER VIA1 ;
        RECT 2.4150 0.5475 2.4900 0.6225 ;
        RECT 1.9575 0.8100 2.0325 0.8850 ;
        RECT 1.1250 0.7950 1.2000 0.8700 ;
        RECT 0.7350 0.3000 0.8100 0.3750 ;
        RECT 0.7275 0.7950 0.8025 0.8700 ;
        LAYER M2 ;
        RECT 2.4000 0.5100 2.5050 0.8850 ;
        RECT 0.7800 0.7800 2.4000 0.8850 ;
        RECT 0.7800 0.3000 0.8850 0.3750 ;
        RECT 0.6900 0.3000 0.7800 0.8850 ;
    END
END OA221_0111


MACRO OA221_1000
    CLASS CORE ;
    FOREIGN OA221_1000 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.6800 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 1.5675 0.1500 1.6425 0.9000 ;
        RECT 1.5375 0.1500 1.5675 0.3825 ;
        RECT 1.5375 0.6675 1.5675 0.9000 ;
        END
    END Z
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.1475 0.8625 1.6125 0.9375 ;
        RECT 1.0725 0.6000 1.1475 0.9375 ;
        RECT 0.7275 0.6000 1.0725 0.6750 ;
        RECT 0.6525 0.4875 0.7275 0.6750 ;
        VIA 0.6900 0.5700 VIA12_square ;
        END
    END C
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.1475 0.2625 1.6125 0.3375 ;
        RECT 1.1475 0.4125 1.2975 0.4875 ;
        RECT 1.0725 0.2625 1.1475 0.4875 ;
        VIA 1.2000 0.4500 VIA12_square ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.8775 0.1125 1.4175 0.1875 ;
        RECT 0.8775 0.4200 0.9675 0.5250 ;
        RECT 0.8025 0.1125 0.8775 0.5250 ;
        VIA 0.8850 0.4725 VIA12_square ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1425 0.4650 0.2475 0.5850 ;
        RECT 0.0675 0.3675 0.1425 0.6825 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.4275 0.1125 0.6075 0.1875 ;
        RECT 0.3525 0.1125 0.4275 0.6600 ;
        RECT 0.0675 0.1125 0.3525 0.1875 ;
        VIA 0.3900 0.5775 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.4250 -0.0750 1.6800 0.0750 ;
        RECT 1.3050 -0.0750 1.4250 0.2475 ;
        RECT 1.0050 -0.0750 1.3050 0.0750 ;
        RECT 0.8850 -0.0750 1.0050 0.1800 ;
        RECT 0.0000 -0.0750 0.8850 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.4250 0.9750 1.6800 1.1250 ;
        RECT 1.3050 0.8325 1.4250 1.1250 ;
        RECT 0.7650 0.9750 1.3050 1.1250 ;
        RECT 0.6600 0.8100 0.7650 1.1250 ;
        RECT 0.1650 0.9750 0.6600 1.1250 ;
        RECT 0.0450 0.8175 0.1650 1.1250 ;
        RECT 0.0000 0.9750 0.0450 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.5450 0.1800 1.6050 0.2400 ;
        RECT 1.5450 0.8100 1.6050 0.8700 ;
        RECT 1.4325 0.4950 1.4925 0.5550 ;
        RECT 1.3350 0.1575 1.3950 0.2175 ;
        RECT 1.3350 0.8325 1.3950 0.8925 ;
        RECT 1.1250 0.1725 1.1850 0.2325 ;
        RECT 1.1250 0.8100 1.1850 0.8700 ;
        RECT 1.0275 0.4950 1.0875 0.5550 ;
        RECT 0.9150 0.1200 0.9750 0.1800 ;
        RECT 0.8100 0.4950 0.8700 0.5550 ;
        RECT 0.7050 0.1800 0.7650 0.2400 ;
        RECT 0.7050 0.8400 0.7650 0.9000 ;
        RECT 0.6000 0.4950 0.6600 0.5550 ;
        RECT 0.4950 0.1575 0.5550 0.2175 ;
        RECT 0.4950 0.8100 0.5550 0.8700 ;
        RECT 0.3900 0.4950 0.4500 0.5550 ;
        RECT 0.2850 0.3075 0.3450 0.3675 ;
        RECT 0.1800 0.4950 0.2400 0.5550 ;
        RECT 0.0750 0.1650 0.1350 0.2250 ;
        RECT 0.0750 0.8325 0.1350 0.8925 ;
        LAYER M1 ;
        RECT 1.4625 0.4650 1.4925 0.5850 ;
        RECT 1.3875 0.4650 1.4625 0.7575 ;
        RECT 1.1925 0.6825 1.3875 0.7575 ;
        RECT 1.0275 0.4125 1.2975 0.6000 ;
        RECT 1.1025 0.1500 1.2075 0.3300 ;
        RECT 1.1175 0.6825 1.1925 0.9000 ;
        RECT 0.8400 0.7875 1.1175 0.9000 ;
        RECT 0.8025 0.2550 1.1025 0.3300 ;
        RECT 0.8100 0.4050 0.9525 0.6975 ;
        RECT 0.6975 0.1500 0.8025 0.3300 ;
        RECT 0.5700 0.4875 0.7275 0.7050 ;
        RECT 0.3825 0.3000 0.6225 0.4125 ;
        RECT 0.1500 0.1500 0.5850 0.2250 ;
        RECT 0.2775 0.7800 0.5850 0.8925 ;
        RECT 0.3300 0.4950 0.4950 0.7050 ;
        RECT 0.2550 0.3000 0.3825 0.3900 ;
        RECT 0.0450 0.1500 0.1500 0.2550 ;
        LAYER VIA1 ;
        RECT 0.8850 0.7875 0.9600 0.8625 ;
        RECT 0.5025 0.3375 0.5775 0.4125 ;
        RECT 0.4275 0.8175 0.5025 0.8925 ;
        LAYER M2 ;
        RECT 0.8400 0.7500 0.9900 0.8925 ;
        RECT 0.5775 0.7500 0.8400 0.8250 ;
        RECT 0.5775 0.2625 0.6075 0.3375 ;
        RECT 0.5025 0.2625 0.5775 0.8925 ;
        RECT 0.3825 0.8175 0.5025 0.8925 ;
    END
END OA221_1000


MACRO OA221_1010
    CLASS CORE ;
    FOREIGN OA221_1010 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.6800 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 1.5675 0.2175 1.6425 0.8325 ;
        RECT 1.5375 0.2175 1.5675 0.3825 ;
        RECT 1.5375 0.6675 1.5675 0.8325 ;
        END
    END Z
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.1475 0.8625 1.6125 0.9375 ;
        RECT 1.0725 0.6000 1.1475 0.9375 ;
        RECT 0.7275 0.6000 1.0725 0.6750 ;
        RECT 0.6525 0.4875 0.7275 0.6750 ;
        VIA 0.6900 0.5700 VIA12_square ;
        END
    END C
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.1475 0.2625 1.6125 0.3375 ;
        RECT 1.1475 0.4125 1.2975 0.4875 ;
        RECT 1.0725 0.2625 1.1475 0.4875 ;
        VIA 1.2000 0.4500 VIA12_square ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.8775 0.1125 1.4175 0.1875 ;
        RECT 0.8775 0.4200 0.9675 0.5250 ;
        RECT 0.8025 0.1125 0.8775 0.5250 ;
        VIA 0.8850 0.4725 VIA12_square ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1425 0.4650 0.2475 0.5850 ;
        RECT 0.0675 0.3675 0.1425 0.6825 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.4275 0.1125 0.6075 0.1875 ;
        RECT 0.3525 0.1125 0.4275 0.6600 ;
        RECT 0.0675 0.1125 0.3525 0.1875 ;
        VIA 0.3900 0.5775 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.4250 -0.0750 1.6800 0.0750 ;
        RECT 1.3050 -0.0750 1.4250 0.3300 ;
        RECT 1.0050 -0.0750 1.3050 0.0750 ;
        RECT 0.8850 -0.0750 1.0050 0.1800 ;
        RECT 0.0000 -0.0750 0.8850 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.4250 0.9750 1.6800 1.1250 ;
        RECT 1.3050 0.8325 1.4250 1.1250 ;
        RECT 0.7650 0.9750 1.3050 1.1250 ;
        RECT 0.6600 0.8100 0.7650 1.1250 ;
        RECT 0.1650 0.9750 0.6600 1.1250 ;
        RECT 0.0450 0.8175 0.1650 1.1250 ;
        RECT 0.0000 0.9750 0.0450 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.5450 0.2700 1.6050 0.3300 ;
        RECT 1.5450 0.7200 1.6050 0.7800 ;
        RECT 1.4325 0.4950 1.4925 0.5550 ;
        RECT 1.3350 0.2400 1.3950 0.3000 ;
        RECT 1.3350 0.8325 1.3950 0.8925 ;
        RECT 1.1250 0.2325 1.1850 0.2925 ;
        RECT 1.1250 0.7725 1.1850 0.8325 ;
        RECT 1.0275 0.4950 1.0875 0.5550 ;
        RECT 0.9150 0.1200 0.9750 0.1800 ;
        RECT 0.8100 0.4950 0.8700 0.5550 ;
        RECT 0.7050 0.2325 0.7650 0.2925 ;
        RECT 0.7050 0.8400 0.7650 0.9000 ;
        RECT 0.6000 0.4950 0.6600 0.5550 ;
        RECT 0.4950 0.1575 0.5550 0.2175 ;
        RECT 0.4950 0.8100 0.5550 0.8700 ;
        RECT 0.3900 0.4950 0.4500 0.5550 ;
        RECT 0.2850 0.3150 0.3450 0.3750 ;
        RECT 0.1800 0.4950 0.2400 0.5550 ;
        RECT 0.0750 0.1650 0.1350 0.2250 ;
        RECT 0.0750 0.8325 0.1350 0.8925 ;
        LAYER M1 ;
        RECT 1.4625 0.4650 1.4925 0.5850 ;
        RECT 1.3875 0.4650 1.4625 0.7575 ;
        RECT 1.1925 0.6825 1.3875 0.7575 ;
        RECT 1.0275 0.4125 1.2975 0.6000 ;
        RECT 1.1175 0.6825 1.1925 0.8925 ;
        RECT 1.0950 0.1950 1.1850 0.3300 ;
        RECT 0.8400 0.7875 1.1175 0.8925 ;
        RECT 0.7950 0.2550 1.0950 0.3300 ;
        RECT 0.8100 0.4050 0.9525 0.6975 ;
        RECT 0.6975 0.2025 0.7950 0.3300 ;
        RECT 0.5700 0.4875 0.7275 0.7050 ;
        RECT 0.3825 0.3000 0.6225 0.4125 ;
        RECT 0.1500 0.1500 0.5850 0.2250 ;
        RECT 0.2775 0.7800 0.5850 0.8925 ;
        RECT 0.3300 0.4950 0.4950 0.7050 ;
        RECT 0.2550 0.3000 0.3825 0.3900 ;
        RECT 0.0450 0.1500 0.1500 0.2550 ;
        LAYER VIA1 ;
        RECT 0.8850 0.7875 0.9600 0.8625 ;
        RECT 0.5025 0.3375 0.5775 0.4125 ;
        RECT 0.4275 0.8175 0.5025 0.8925 ;
        LAYER M2 ;
        RECT 0.8400 0.7500 0.9900 0.8925 ;
        RECT 0.5775 0.7500 0.8400 0.8250 ;
        RECT 0.5775 0.2625 0.6075 0.3375 ;
        RECT 0.5025 0.2625 0.5775 0.8925 ;
        RECT 0.3825 0.8175 0.5025 0.8925 ;
    END
END OA221_1010


MACRO OA222_0011
    CLASS CORE ;
    FOREIGN OA222_0011 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.1000 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 1.9875 0.3075 2.0625 0.7425 ;
        RECT 1.8225 0.3075 1.9875 0.3825 ;
        RECT 1.8225 0.6675 1.9875 0.7425 ;
        RECT 1.7475 0.2175 1.8225 0.3825 ;
        RECT 1.7475 0.6675 1.8225 0.8550 ;
        END
    END Z
    PIN C2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.0725 0.5625 1.5375 0.6375 ;
        VIA 1.2225 0.6000 VIA12_square ;
        END
    END C2
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.2750 0.4125 1.8225 0.4875 ;
        VIA 1.4850 0.4500 VIA12_square ;
        END
    END C1
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.6075 0.5550 0.6375 0.7050 ;
        RECT 0.5325 0.5550 0.6075 0.9375 ;
        RECT 0.0675 0.8625 0.5325 0.9375 ;
        VIA 0.5850 0.6300 VIA12_square ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.9525 0.1125 1.2750 0.1875 ;
        RECT 0.8775 0.1125 0.9525 0.7050 ;
        RECT 0.7200 0.1125 0.8775 0.1875 ;
        VIA 0.9150 0.5925 VIA12_square ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1425 0.4650 0.2475 0.5850 ;
        RECT 0.0675 0.3675 0.1425 0.6825 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.4275 0.1125 0.6000 0.1875 ;
        RECT 0.3525 0.1125 0.4275 0.7125 ;
        RECT 0.0600 0.1125 0.3525 0.1875 ;
        VIA 0.3900 0.6300 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 2.0550 -0.0750 2.1000 0.0750 ;
        RECT 1.9350 -0.0750 2.0550 0.2175 ;
        RECT 1.6350 -0.0750 1.9350 0.0750 ;
        RECT 1.5150 -0.0750 1.6350 0.1800 ;
        RECT 1.2150 -0.0750 1.5150 0.0750 ;
        RECT 1.0950 -0.0750 1.2150 0.2175 ;
        RECT 0.0000 -0.0750 1.0950 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 2.0550 0.9750 2.1000 1.1250 ;
        RECT 1.9350 0.8175 2.0550 1.1250 ;
        RECT 1.6350 0.9750 1.9350 1.1250 ;
        RECT 1.5150 0.8700 1.6350 1.1250 ;
        RECT 1.0200 0.9750 1.5150 1.1250 ;
        RECT 0.9150 0.7875 1.0200 1.1250 ;
        RECT 0.1650 0.9750 0.9150 1.1250 ;
        RECT 0.0450 0.7875 0.1650 1.1250 ;
        RECT 0.0000 0.9750 0.0450 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.9650 0.1575 2.0250 0.2175 ;
        RECT 1.9650 0.8325 2.0250 0.8925 ;
        RECT 1.8525 0.4950 1.9125 0.5550 ;
        RECT 1.7550 0.2775 1.8150 0.3375 ;
        RECT 1.7550 0.7650 1.8150 0.8250 ;
        RECT 1.6500 0.4950 1.7100 0.5550 ;
        RECT 1.5450 0.1200 1.6050 0.1800 ;
        RECT 1.5450 0.8700 1.6050 0.9300 ;
        RECT 1.4400 0.5025 1.5000 0.5625 ;
        RECT 1.3350 0.1725 1.3950 0.2325 ;
        RECT 1.2225 0.5025 1.2825 0.5625 ;
        RECT 1.1250 0.1575 1.1850 0.2175 ;
        RECT 1.1250 0.8100 1.1850 0.8700 ;
        RECT 0.9150 0.1800 0.9750 0.2400 ;
        RECT 0.9150 0.8325 0.9750 0.8925 ;
        RECT 0.8100 0.5025 0.8700 0.5625 ;
        RECT 0.7050 0.3300 0.7650 0.3900 ;
        RECT 0.6000 0.5025 0.6600 0.5625 ;
        RECT 0.4950 0.1575 0.5550 0.2175 ;
        RECT 0.4950 0.8250 0.5550 0.8850 ;
        RECT 0.3900 0.4950 0.4500 0.5550 ;
        RECT 0.2850 0.3225 0.3450 0.3825 ;
        RECT 0.1800 0.4950 0.2400 0.5550 ;
        RECT 0.0750 0.1725 0.1350 0.2325 ;
        RECT 0.0750 0.8175 0.1350 0.8775 ;
        LAYER M1 ;
        RECT 1.6725 0.4650 1.9125 0.5850 ;
        RECT 1.5975 0.4650 1.6725 0.7950 ;
        RECT 1.4400 0.7200 1.5975 0.7950 ;
        RECT 1.4400 0.3675 1.5225 0.6450 ;
        RECT 1.3575 0.4500 1.4400 0.6450 ;
        RECT 1.3650 0.7200 1.4400 0.9000 ;
        RECT 1.3650 0.1500 1.4250 0.2550 ;
        RECT 1.2900 0.1500 1.3650 0.3675 ;
        RECT 1.0950 0.7950 1.3650 0.9000 ;
        RECT 1.1400 0.2925 1.2900 0.3675 ;
        RECT 1.2000 0.4725 1.2825 0.7050 ;
        RECT 1.0500 0.4950 1.2000 0.7050 ;
        RECT 1.0650 0.2925 1.1400 0.4200 ;
        RECT 0.8100 0.3450 1.0650 0.4200 ;
        RECT 0.8850 0.1500 0.9900 0.2700 ;
        RECT 0.7800 0.4950 0.9750 0.7050 ;
        RECT 0.1575 0.1500 0.8850 0.2250 ;
        RECT 0.6600 0.7800 0.8400 0.8925 ;
        RECT 0.7050 0.3000 0.8100 0.4200 ;
        RECT 0.5325 0.4950 0.6975 0.7050 ;
        RECT 0.3750 0.8175 0.6600 0.8925 ;
        RECT 0.5100 0.3000 0.6300 0.4200 ;
        RECT 0.2550 0.3000 0.5100 0.3900 ;
        RECT 0.3300 0.4650 0.4500 0.7425 ;
        RECT 0.0525 0.1500 0.1575 0.2550 ;
        LAYER VIA1 ;
        RECT 1.1400 0.8100 1.2150 0.8850 ;
        RECT 0.7125 0.7875 0.7875 0.8625 ;
        RECT 0.5100 0.3075 0.5850 0.3825 ;
        LAYER M2 ;
        RECT 1.1025 0.7950 1.2525 0.9000 ;
        RECT 0.8025 0.8250 1.1025 0.9000 ;
        RECT 0.7275 0.2625 0.8025 0.9000 ;
        RECT 0.6075 0.2625 0.7275 0.3375 ;
        RECT 0.6975 0.7500 0.7275 0.9000 ;
        RECT 0.5025 0.2625 0.6075 0.4275 ;
    END
END OA222_0011


MACRO OA222_0111
    CLASS CORE ;
    FOREIGN OA222_0111 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.7800 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 3.0975 0.2400 3.4125 0.7500 ;
        VIA 3.2550 0.3225 VIA12_slot ;
        VIA 3.2550 0.6675 VIA12_slot ;
        END
    END Z
    PIN C2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 2.3775 0.2625 2.4525 0.6075 ;
        RECT 1.9050 0.2625 2.3775 0.3375 ;
        VIA 2.4150 0.5250 VIA12_square ;
        END
    END C2
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.6650 0.5625 2.1375 0.6375 ;
        VIA 2.0400 0.6000 VIA12_square ;
        END
    END C1
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.4025 0.4125 1.8750 0.4875 ;
        RECT 1.3275 0.4125 1.4025 0.6000 ;
        VIA 1.3650 0.5175 VIA12_square ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.0125 0.1125 1.0875 0.6675 ;
        RECT 0.5475 0.1125 1.0125 0.1875 ;
        VIA 1.0500 0.5700 VIA12_square ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.7875 0.4725 0.8925 0.7200 ;
        RECT 0.2400 0.6450 0.7875 0.7200 ;
        RECT 0.1425 0.4650 0.2400 0.7200 ;
        RECT 0.0675 0.3675 0.1425 0.7200 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.5325 0.3975 0.6075 0.7875 ;
        RECT 0.0675 0.7125 0.5325 0.7875 ;
        VIA 0.5700 0.5175 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 3.7125 -0.0750 3.7800 0.0750 ;
        RECT 3.6375 -0.0750 3.7125 0.3150 ;
        RECT 3.3150 -0.0750 3.6375 0.0750 ;
        RECT 3.1950 -0.0750 3.3150 0.1950 ;
        RECT 2.8950 -0.0750 3.1950 0.0750 ;
        RECT 2.7750 -0.0750 2.8950 0.2475 ;
        RECT 2.4750 -0.0750 2.7750 0.0750 ;
        RECT 2.3550 -0.0750 2.4750 0.2325 ;
        RECT 2.0550 -0.0750 2.3550 0.0750 ;
        RECT 1.9500 -0.0750 2.0550 0.2475 ;
        RECT 0.0000 -0.0750 1.9500 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 3.7125 0.9750 3.7800 1.1250 ;
        RECT 3.6375 0.6375 3.7125 1.1250 ;
        RECT 3.3075 0.9750 3.6375 1.1250 ;
        RECT 3.2025 0.8025 3.3075 1.1250 ;
        RECT 2.8725 0.9750 3.2025 1.1250 ;
        RECT 2.7975 0.6750 2.8725 1.1250 ;
        RECT 2.0550 0.9750 2.7975 1.1250 ;
        RECT 1.9350 0.8025 2.0550 1.1250 ;
        RECT 1.8450 0.9750 1.9350 1.1250 ;
        RECT 1.7250 0.8025 1.8450 1.1250 ;
        RECT 1.0200 0.9750 1.7250 1.1250 ;
        RECT 0.9150 0.7950 1.0200 1.1250 ;
        RECT 0.1575 0.9750 0.9150 1.1250 ;
        RECT 0.0525 0.8025 0.1575 1.1250 ;
        RECT 0.0000 0.9750 0.0525 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 3.6450 0.2250 3.7050 0.2850 ;
        RECT 3.6450 0.6675 3.7050 0.7275 ;
        RECT 3.6450 0.8325 3.7050 0.8925 ;
        RECT 3.5400 0.4650 3.6000 0.5250 ;
        RECT 3.4350 0.2250 3.4950 0.2850 ;
        RECT 3.4350 0.7575 3.4950 0.8175 ;
        RECT 3.3300 0.4650 3.3900 0.5250 ;
        RECT 3.2250 0.1275 3.2850 0.1875 ;
        RECT 3.2250 0.8325 3.2850 0.8925 ;
        RECT 3.1200 0.4650 3.1800 0.5250 ;
        RECT 3.0150 0.2250 3.0750 0.2850 ;
        RECT 3.0150 0.7575 3.0750 0.8175 ;
        RECT 2.9100 0.4650 2.9700 0.5250 ;
        RECT 2.8050 0.1650 2.8650 0.2250 ;
        RECT 2.8050 0.7050 2.8650 0.7650 ;
        RECT 2.8050 0.8700 2.8650 0.9300 ;
        RECT 2.7000 0.4875 2.7600 0.5475 ;
        RECT 2.5950 0.3150 2.6550 0.3750 ;
        RECT 2.4900 0.4950 2.5500 0.5550 ;
        RECT 2.3850 0.1575 2.4450 0.2175 ;
        RECT 2.3850 0.8175 2.4450 0.8775 ;
        RECT 2.2800 0.4950 2.3400 0.5550 ;
        RECT 2.1750 0.3150 2.2350 0.3750 ;
        RECT 2.0700 0.4950 2.1300 0.5550 ;
        RECT 1.9650 0.1575 2.0250 0.2175 ;
        RECT 1.9650 0.8175 2.0250 0.8775 ;
        RECT 1.7550 0.1575 1.8150 0.2175 ;
        RECT 1.7550 0.8175 1.8150 0.8775 ;
        RECT 1.6500 0.4950 1.7100 0.5550 ;
        RECT 1.5450 0.3225 1.6050 0.3825 ;
        RECT 1.4400 0.4950 1.5000 0.5550 ;
        RECT 1.3350 0.1575 1.3950 0.2175 ;
        RECT 1.3350 0.8100 1.3950 0.8700 ;
        RECT 1.2300 0.4950 1.2900 0.5550 ;
        RECT 1.1250 0.3225 1.1850 0.3825 ;
        RECT 1.0200 0.4950 1.0800 0.5550 ;
        RECT 0.9150 0.1575 0.9750 0.2175 ;
        RECT 0.9150 0.8250 0.9750 0.8850 ;
        RECT 0.8100 0.4950 0.8700 0.5550 ;
        RECT 0.7050 0.3150 0.7650 0.3750 ;
        RECT 0.6000 0.4950 0.6600 0.5550 ;
        RECT 0.4950 0.1575 0.5550 0.2175 ;
        RECT 0.4950 0.8175 0.5550 0.8775 ;
        RECT 0.3900 0.4950 0.4500 0.5550 ;
        RECT 0.2850 0.3150 0.3450 0.3750 ;
        RECT 0.1800 0.4950 0.2400 0.5550 ;
        RECT 0.0750 0.1725 0.1350 0.2325 ;
        RECT 0.0750 0.8325 0.1350 0.8925 ;
        LAYER M1 ;
        RECT 2.9100 0.4425 3.6300 0.5475 ;
        RECT 3.4125 0.1950 3.5175 0.3675 ;
        RECT 3.4275 0.6225 3.5025 0.8700 ;
        RECT 3.0825 0.6225 3.4275 0.7125 ;
        RECT 3.0975 0.2775 3.4125 0.3675 ;
        RECT 2.9925 0.1950 3.0975 0.3675 ;
        RECT 3.0075 0.6225 3.0825 0.8700 ;
        RECT 2.8350 0.3750 2.9100 0.5475 ;
        RECT 2.7225 0.4575 2.7600 0.5775 ;
        RECT 2.6475 0.4575 2.7225 0.7275 ;
        RECT 2.2125 0.3075 2.6850 0.3825 ;
        RECT 2.1600 0.6525 2.6475 0.7275 ;
        RECT 2.2425 0.8025 2.5875 0.9000 ;
        RECT 2.2500 0.4725 2.5725 0.5775 ;
        RECT 2.1375 0.3075 2.2125 0.3975 ;
        RECT 2.0550 0.4875 2.1600 0.7275 ;
        RECT 1.8750 0.3225 2.1375 0.3975 ;
        RECT 1.9575 0.4875 2.0550 0.6600 ;
        RECT 1.8075 0.3150 1.8750 0.3975 ;
        RECT 0.1575 0.1500 1.8450 0.2250 ;
        RECT 1.0725 0.3150 1.8075 0.3900 ;
        RECT 1.6275 0.4725 1.7325 0.7200 ;
        RECT 1.1025 0.6450 1.6275 0.7200 ;
        RECT 1.2000 0.4650 1.5300 0.5700 ;
        RECT 1.2075 0.7950 1.5075 0.9000 ;
        RECT 0.9975 0.4650 1.1025 0.7200 ;
        RECT 0.2475 0.3075 0.8475 0.3900 ;
        RECT 0.4650 0.7950 0.8400 0.9000 ;
        RECT 0.3600 0.4650 0.6900 0.5700 ;
        RECT 0.0525 0.1500 0.1575 0.2550 ;
        LAYER VIA1 ;
        RECT 2.8350 0.4275 2.9100 0.5025 ;
        RECT 2.3775 0.8100 2.4525 0.8850 ;
        RECT 1.3275 0.8025 1.4025 0.8775 ;
        RECT 0.7275 0.3150 0.8025 0.3900 ;
        RECT 0.7275 0.8100 0.8025 0.8850 ;
        LAYER M2 ;
        RECT 2.8200 0.3900 2.9250 0.8850 ;
        RECT 0.8400 0.7950 2.8200 0.8850 ;
        RECT 0.7875 0.3075 0.8475 0.3900 ;
        RECT 0.7875 0.7950 0.8400 0.9000 ;
        RECT 0.6825 0.3075 0.7875 0.9000 ;
    END
END OA222_0111


MACRO OA222_1000
    CLASS CORE ;
    FOREIGN OA222_1000 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.8900 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 1.7775 0.1500 1.8525 0.9000 ;
        RECT 1.7475 0.1500 1.7775 0.3825 ;
        RECT 1.7475 0.6675 1.7775 0.9000 ;
        END
    END Z
    PIN C2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.0725 0.5625 1.5375 0.6375 ;
        VIA 1.2225 0.6000 VIA12_square ;
        END
    END C2
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.2750 0.4125 1.7400 0.4875 ;
        VIA 1.4850 0.4500 VIA12_square ;
        END
    END C1
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.6075 0.5550 0.6375 0.7050 ;
        RECT 0.5325 0.5550 0.6075 0.9375 ;
        RECT 0.0675 0.8625 0.5325 0.9375 ;
        VIA 0.5850 0.6300 VIA12_square ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.9525 0.1125 1.2750 0.1875 ;
        RECT 0.8775 0.1125 0.9525 0.7050 ;
        RECT 0.7200 0.1125 0.8775 0.1875 ;
        VIA 0.9150 0.5925 VIA12_square ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1425 0.4650 0.2475 0.5850 ;
        RECT 0.0675 0.3675 0.1425 0.6825 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.4275 0.1125 0.6000 0.1875 ;
        RECT 0.3525 0.1125 0.4275 0.7125 ;
        RECT 0.0600 0.1125 0.3525 0.1875 ;
        VIA 0.3900 0.6300 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.6350 -0.0750 1.8900 0.0750 ;
        RECT 1.5150 -0.0750 1.6350 0.1800 ;
        RECT 1.2150 -0.0750 1.5150 0.0750 ;
        RECT 1.0950 -0.0750 1.2150 0.2175 ;
        RECT 0.0000 -0.0750 1.0950 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.6350 0.9750 1.8900 1.1250 ;
        RECT 1.5150 0.8700 1.6350 1.1250 ;
        RECT 1.0200 0.9750 1.5150 1.1250 ;
        RECT 0.9150 0.7875 1.0200 1.1250 ;
        RECT 0.1650 0.9750 0.9150 1.1250 ;
        RECT 0.0450 0.7875 0.1650 1.1250 ;
        RECT 0.0000 0.9750 0.0450 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.7550 0.1800 1.8150 0.2400 ;
        RECT 1.7550 0.8100 1.8150 0.8700 ;
        RECT 1.6425 0.4950 1.7025 0.5550 ;
        RECT 1.5450 0.1200 1.6050 0.1800 ;
        RECT 1.5450 0.8700 1.6050 0.9300 ;
        RECT 1.4400 0.5025 1.5000 0.5625 ;
        RECT 1.3350 0.1725 1.3950 0.2325 ;
        RECT 1.2225 0.5025 1.2825 0.5625 ;
        RECT 1.1250 0.1575 1.1850 0.2175 ;
        RECT 1.1250 0.8100 1.1850 0.8700 ;
        RECT 0.9150 0.1800 0.9750 0.2400 ;
        RECT 0.9150 0.8325 0.9750 0.8925 ;
        RECT 0.8100 0.5025 0.8700 0.5625 ;
        RECT 0.7050 0.3300 0.7650 0.3900 ;
        RECT 0.6000 0.5025 0.6600 0.5625 ;
        RECT 0.4950 0.1650 0.5550 0.2250 ;
        RECT 0.4950 0.8250 0.5550 0.8850 ;
        RECT 0.3900 0.4950 0.4500 0.5550 ;
        RECT 0.2850 0.3225 0.3450 0.3825 ;
        RECT 0.1800 0.4950 0.2400 0.5550 ;
        RECT 0.0750 0.1800 0.1350 0.2400 ;
        RECT 0.0750 0.8175 0.1350 0.8775 ;
        LAYER M1 ;
        RECT 1.6725 0.4650 1.7025 0.5850 ;
        RECT 1.5975 0.4650 1.6725 0.7950 ;
        RECT 1.4400 0.7200 1.5975 0.7950 ;
        RECT 1.4400 0.3675 1.5225 0.6450 ;
        RECT 1.3575 0.4500 1.4400 0.6450 ;
        RECT 1.3650 0.7200 1.4400 0.9000 ;
        RECT 1.3650 0.1500 1.4250 0.2550 ;
        RECT 1.2900 0.1500 1.3650 0.3675 ;
        RECT 1.0950 0.7950 1.3650 0.9000 ;
        RECT 1.1400 0.2925 1.2900 0.3675 ;
        RECT 1.2000 0.4725 1.2825 0.7050 ;
        RECT 1.0500 0.4950 1.2000 0.7050 ;
        RECT 1.0650 0.2925 1.1400 0.4200 ;
        RECT 0.8100 0.3450 1.0650 0.4200 ;
        RECT 0.8850 0.1500 0.9900 0.2700 ;
        RECT 0.7800 0.4950 0.9750 0.7050 ;
        RECT 0.1575 0.1500 0.8850 0.2250 ;
        RECT 0.6600 0.7800 0.8400 0.8925 ;
        RECT 0.7050 0.3000 0.8100 0.4200 ;
        RECT 0.5325 0.4950 0.6975 0.7050 ;
        RECT 0.3750 0.8175 0.6600 0.8925 ;
        RECT 0.5100 0.3000 0.6300 0.4200 ;
        RECT 0.2550 0.3000 0.5100 0.3900 ;
        RECT 0.3300 0.4650 0.4500 0.7425 ;
        RECT 0.0525 0.1500 0.1575 0.2625 ;
        LAYER VIA1 ;
        RECT 1.1400 0.8100 1.2150 0.8850 ;
        RECT 0.7125 0.7875 0.7875 0.8625 ;
        RECT 0.5100 0.3075 0.5850 0.3825 ;
        LAYER M2 ;
        RECT 1.1025 0.7950 1.2525 0.9000 ;
        RECT 0.8025 0.8250 1.1025 0.9000 ;
        RECT 0.7275 0.2625 0.8025 0.9000 ;
        RECT 0.6075 0.2625 0.7275 0.3375 ;
        RECT 0.6975 0.7500 0.7275 0.9000 ;
        RECT 0.5025 0.2625 0.6075 0.4275 ;
    END
END OA222_1000


MACRO OA222_1010
    CLASS CORE ;
    FOREIGN OA222_1010 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.8900 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 1.7775 0.2175 1.8525 0.8325 ;
        RECT 1.7475 0.2175 1.7775 0.3825 ;
        RECT 1.7475 0.6675 1.7775 0.8325 ;
        END
    END Z
    PIN C2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.0725 0.5625 1.5375 0.6375 ;
        VIA 1.2225 0.6000 VIA12_square ;
        END
    END C2
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.2750 0.4125 1.7400 0.4875 ;
        VIA 1.4850 0.4500 VIA12_square ;
        END
    END C1
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.6075 0.5550 0.6375 0.7050 ;
        RECT 0.5325 0.5550 0.6075 0.9375 ;
        RECT 0.0675 0.8625 0.5325 0.9375 ;
        VIA 0.5850 0.6300 VIA12_square ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.9525 0.1125 1.2750 0.1875 ;
        RECT 0.8775 0.1125 0.9525 0.7050 ;
        RECT 0.7200 0.1125 0.8775 0.1875 ;
        VIA 0.9150 0.5925 VIA12_square ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1425 0.4650 0.2475 0.5850 ;
        RECT 0.0675 0.3675 0.1425 0.6825 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.4275 0.1125 0.6000 0.1875 ;
        RECT 0.3525 0.1125 0.4275 0.7125 ;
        RECT 0.0600 0.1125 0.3525 0.1875 ;
        VIA 0.3900 0.6300 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.6350 -0.0750 1.8900 0.0750 ;
        RECT 1.5150 -0.0750 1.6350 0.1800 ;
        RECT 1.2150 -0.0750 1.5150 0.0750 ;
        RECT 1.0950 -0.0750 1.2150 0.2175 ;
        RECT 0.0000 -0.0750 1.0950 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.6350 0.9750 1.8900 1.1250 ;
        RECT 1.5150 0.8700 1.6350 1.1250 ;
        RECT 1.0200 0.9750 1.5150 1.1250 ;
        RECT 0.9150 0.7875 1.0200 1.1250 ;
        RECT 0.1650 0.9750 0.9150 1.1250 ;
        RECT 0.0450 0.7875 0.1650 1.1250 ;
        RECT 0.0000 0.9750 0.0450 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.7550 0.2700 1.8150 0.3300 ;
        RECT 1.7550 0.7200 1.8150 0.7800 ;
        RECT 1.6425 0.4950 1.7025 0.5550 ;
        RECT 1.5450 0.1200 1.6050 0.1800 ;
        RECT 1.5450 0.8700 1.6050 0.9300 ;
        RECT 1.4400 0.5025 1.5000 0.5625 ;
        RECT 1.3350 0.1725 1.3950 0.2325 ;
        RECT 1.2225 0.5025 1.2825 0.5625 ;
        RECT 1.1250 0.1575 1.1850 0.2175 ;
        RECT 1.1250 0.8100 1.1850 0.8700 ;
        RECT 0.9150 0.1800 0.9750 0.2400 ;
        RECT 0.9150 0.8325 0.9750 0.8925 ;
        RECT 0.8100 0.5025 0.8700 0.5625 ;
        RECT 0.7050 0.3300 0.7650 0.3900 ;
        RECT 0.6000 0.5025 0.6600 0.5625 ;
        RECT 0.4950 0.1575 0.5550 0.2175 ;
        RECT 0.4950 0.8250 0.5550 0.8850 ;
        RECT 0.3900 0.4950 0.4500 0.5550 ;
        RECT 0.2850 0.3225 0.3450 0.3825 ;
        RECT 0.1800 0.4950 0.2400 0.5550 ;
        RECT 0.0750 0.1725 0.1350 0.2325 ;
        RECT 0.0750 0.8175 0.1350 0.8775 ;
        LAYER M1 ;
        RECT 1.6725 0.4650 1.7025 0.5850 ;
        RECT 1.5975 0.4650 1.6725 0.7950 ;
        RECT 1.4400 0.7200 1.5975 0.7950 ;
        RECT 1.4400 0.3675 1.5225 0.6450 ;
        RECT 1.3575 0.4500 1.4400 0.6450 ;
        RECT 1.3650 0.7200 1.4400 0.9000 ;
        RECT 1.3650 0.1500 1.4250 0.2550 ;
        RECT 1.2900 0.1500 1.3650 0.3675 ;
        RECT 1.0950 0.7950 1.3650 0.9000 ;
        RECT 1.1400 0.2925 1.2900 0.3675 ;
        RECT 1.2000 0.4725 1.2825 0.7050 ;
        RECT 1.0500 0.4950 1.2000 0.7050 ;
        RECT 1.0650 0.2925 1.1400 0.4200 ;
        RECT 0.8100 0.3450 1.0650 0.4200 ;
        RECT 0.8850 0.1500 0.9900 0.2700 ;
        RECT 0.7800 0.4950 0.9750 0.7050 ;
        RECT 0.1575 0.1500 0.8850 0.2250 ;
        RECT 0.6600 0.7800 0.8400 0.8925 ;
        RECT 0.7050 0.3000 0.8100 0.4200 ;
        RECT 0.5325 0.4950 0.6975 0.7050 ;
        RECT 0.3750 0.8175 0.6600 0.8925 ;
        RECT 0.5100 0.3000 0.6300 0.4200 ;
        RECT 0.2550 0.3000 0.5100 0.3900 ;
        RECT 0.3300 0.4650 0.4500 0.7425 ;
        RECT 0.0525 0.1500 0.1575 0.2550 ;
        LAYER VIA1 ;
        RECT 1.1400 0.8100 1.2150 0.8850 ;
        RECT 0.7125 0.7875 0.7875 0.8625 ;
        RECT 0.5100 0.3075 0.5850 0.3825 ;
        LAYER M2 ;
        RECT 1.1025 0.7950 1.2525 0.9000 ;
        RECT 0.8025 0.8250 1.1025 0.9000 ;
        RECT 0.7275 0.2625 0.8025 0.9000 ;
        RECT 0.6075 0.2625 0.7275 0.3375 ;
        RECT 0.6975 0.7500 0.7275 0.9000 ;
        RECT 0.5025 0.2625 0.6075 0.4275 ;
    END
END OA222_1010


MACRO OA22_0011
    CLASS CORE ;
    FOREIGN OA22_0011 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.6800 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 1.5675 0.3075 1.6425 0.7425 ;
        RECT 1.4025 0.3075 1.5675 0.3825 ;
        RECT 1.4025 0.6675 1.5675 0.7425 ;
        RECT 1.3275 0.2175 1.4025 0.3825 ;
        RECT 1.3275 0.6675 1.4025 0.8550 ;
        END
    END Z
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.8775 0.4125 1.3425 0.4875 ;
        VIA 0.9900 0.4500 VIA12_square ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.7575 0.1125 1.2075 0.1875 ;
        RECT 0.6525 0.1125 0.7575 0.5700 ;
        VIA 0.7050 0.4875 VIA12_square ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1425 0.5100 0.2700 0.6150 ;
        RECT 0.0675 0.3675 0.1425 0.6825 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.5775 0.7125 1.0950 0.7875 ;
        RECT 0.5025 0.5550 0.5775 0.7875 ;
        VIA 0.5400 0.6750 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.6350 -0.0750 1.6800 0.0750 ;
        RECT 1.5150 -0.0750 1.6350 0.2175 ;
        RECT 1.2150 -0.0750 1.5150 0.0750 ;
        RECT 1.0950 -0.0750 1.2150 0.2475 ;
        RECT 0.7950 -0.0750 1.0950 0.0750 ;
        RECT 0.6750 -0.0750 0.7950 0.1800 ;
        RECT 0.0000 -0.0750 0.6750 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.6350 0.9750 1.6800 1.1250 ;
        RECT 1.5150 0.8175 1.6350 1.1250 ;
        RECT 1.2150 0.9750 1.5150 1.1250 ;
        RECT 1.0950 0.8325 1.2150 1.1250 ;
        RECT 1.0050 0.9750 1.0950 1.1250 ;
        RECT 0.8850 0.8325 1.0050 1.1250 ;
        RECT 0.1650 0.9750 0.8850 1.1250 ;
        RECT 0.0450 0.8025 0.1650 1.1250 ;
        RECT 0.0000 0.9750 0.0450 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.5450 0.1575 1.6050 0.2175 ;
        RECT 1.5450 0.8325 1.6050 0.8925 ;
        RECT 1.4325 0.4950 1.4925 0.5550 ;
        RECT 1.3350 0.2775 1.3950 0.3375 ;
        RECT 1.3350 0.7650 1.3950 0.8250 ;
        RECT 1.2300 0.4950 1.2900 0.5550 ;
        RECT 1.1250 0.1575 1.1850 0.2175 ;
        RECT 1.1250 0.8325 1.1850 0.8925 ;
        RECT 0.9150 0.2325 0.9750 0.2925 ;
        RECT 0.9150 0.8325 0.9750 0.8925 ;
        RECT 0.8175 0.4950 0.8775 0.5550 ;
        RECT 0.7050 0.1200 0.7650 0.1800 ;
        RECT 0.6000 0.4950 0.6600 0.5550 ;
        RECT 0.4950 0.1575 0.5550 0.2175 ;
        RECT 0.4950 0.7950 0.5550 0.8550 ;
        RECT 0.3825 0.5400 0.4425 0.6000 ;
        RECT 0.2850 0.3375 0.3450 0.3975 ;
        RECT 0.1800 0.5100 0.2400 0.5700 ;
        RECT 0.0750 0.8325 0.1350 0.8925 ;
        RECT 0.0750 0.1650 0.1350 0.2250 ;
        LAYER M1 ;
        RECT 1.2525 0.4650 1.4925 0.5850 ;
        RECT 1.1775 0.4650 1.2525 0.7575 ;
        RECT 0.8100 0.6825 1.1775 0.7575 ;
        RECT 0.8175 0.4125 1.0875 0.6000 ;
        RECT 0.8850 0.1950 0.9750 0.3300 ;
        RECT 0.6000 0.2550 0.8850 0.3300 ;
        RECT 0.7350 0.6825 0.8100 0.8625 ;
        RECT 0.6675 0.4050 0.7425 0.5775 ;
        RECT 0.3075 0.7875 0.7350 0.8625 ;
        RECT 0.5475 0.4050 0.6675 0.5625 ;
        RECT 0.4725 0.6375 0.6225 0.7125 ;
        RECT 0.5250 0.1500 0.6000 0.3300 ;
        RECT 0.1500 0.1500 0.5250 0.2250 ;
        RECT 0.3525 0.5400 0.4725 0.7125 ;
        RECT 0.3450 0.3000 0.4500 0.4650 ;
        RECT 0.2175 0.3000 0.3450 0.4350 ;
        RECT 0.0450 0.1500 0.1500 0.2550 ;
        LAYER VIA1 ;
        RECT 0.3525 0.3450 0.4275 0.4200 ;
        RECT 0.3525 0.7875 0.4275 0.8625 ;
        LAYER M2 ;
        RECT 0.4275 0.8625 0.4575 0.9375 ;
        RECT 0.3525 0.3000 0.4275 0.9375 ;
    END
END OA22_0011


MACRO OA22_0111
    CLASS CORE ;
    FOREIGN OA22_0111 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.9400 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 2.2575 0.2400 2.5725 0.7500 ;
        VIA 2.4150 0.3225 VIA12_slot ;
        VIA 2.4150 0.6675 VIA12_slot ;
        END
    END Z
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.1175 0.1125 1.1925 0.6675 ;
        RECT 0.6525 0.1125 1.1175 0.1875 ;
        VIA 1.1550 0.5775 VIA12_square ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.6125 0.2625 2.0850 0.3375 ;
        RECT 1.5375 0.2625 1.6125 0.6075 ;
        VIA 1.5750 0.5250 VIA12_square ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.7875 0.4725 0.8925 0.7050 ;
        RECT 0.2400 0.6300 0.7875 0.7050 ;
        RECT 0.1425 0.4650 0.2400 0.7050 ;
        RECT 0.0675 0.3675 0.1425 0.7050 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.4950 0.3975 0.6000 0.7875 ;
        RECT 0.0675 0.7125 0.4950 0.7875 ;
        VIA 0.5475 0.5025 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 2.8725 -0.0750 2.9400 0.0750 ;
        RECT 2.7975 -0.0750 2.8725 0.3150 ;
        RECT 2.4750 -0.0750 2.7975 0.0750 ;
        RECT 2.3550 -0.0750 2.4750 0.1950 ;
        RECT 2.0325 -0.0750 2.3550 0.0750 ;
        RECT 1.9575 -0.0750 2.0325 0.2925 ;
        RECT 1.6350 -0.0750 1.9575 0.0750 ;
        RECT 1.5150 -0.0750 1.6350 0.2400 ;
        RECT 1.2075 -0.0750 1.5150 0.0750 ;
        RECT 1.1025 -0.0750 1.2075 0.2400 ;
        RECT 0.0000 -0.0750 1.1025 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 2.8725 0.9750 2.9400 1.1250 ;
        RECT 2.7975 0.6375 2.8725 1.1250 ;
        RECT 2.4525 0.9750 2.7975 1.1250 ;
        RECT 2.3775 0.8175 2.4525 1.1250 ;
        RECT 2.0550 0.9750 2.3775 1.1250 ;
        RECT 1.9350 0.8025 2.0550 1.1250 ;
        RECT 1.2150 0.9750 1.9350 1.1250 ;
        RECT 1.0950 0.8025 1.2150 1.1250 ;
        RECT 1.0200 0.9750 1.0950 1.1250 ;
        RECT 0.9150 0.7950 1.0200 1.1250 ;
        RECT 0.1575 0.9750 0.9150 1.1250 ;
        RECT 0.0525 0.8025 0.1575 1.1250 ;
        RECT 0.0000 0.9750 0.0525 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 2.8050 0.2250 2.8650 0.2850 ;
        RECT 2.8050 0.6675 2.8650 0.7275 ;
        RECT 2.8050 0.8325 2.8650 0.8925 ;
        RECT 2.7000 0.4650 2.7600 0.5250 ;
        RECT 2.5950 0.2250 2.6550 0.2850 ;
        RECT 2.5950 0.7575 2.6550 0.8175 ;
        RECT 2.4900 0.4650 2.5500 0.5250 ;
        RECT 2.3850 0.1275 2.4450 0.1875 ;
        RECT 2.3850 0.8475 2.4450 0.9075 ;
        RECT 2.2800 0.4650 2.3400 0.5250 ;
        RECT 2.1750 0.2250 2.2350 0.2850 ;
        RECT 2.1750 0.7575 2.2350 0.8175 ;
        RECT 2.0700 0.4650 2.1300 0.5250 ;
        RECT 1.9650 0.2025 2.0250 0.2625 ;
        RECT 1.9650 0.8250 2.0250 0.8850 ;
        RECT 1.8600 0.4950 1.9200 0.5550 ;
        RECT 1.7550 0.3225 1.8150 0.3825 ;
        RECT 1.6500 0.4950 1.7100 0.5550 ;
        RECT 1.5450 0.1575 1.6050 0.2175 ;
        RECT 1.5450 0.8175 1.6050 0.8775 ;
        RECT 1.4400 0.4950 1.5000 0.5550 ;
        RECT 1.3350 0.3225 1.3950 0.3825 ;
        RECT 1.2300 0.4950 1.2900 0.5550 ;
        RECT 1.1250 0.1575 1.1850 0.2175 ;
        RECT 1.1250 0.8175 1.1850 0.8775 ;
        RECT 0.9150 0.2400 0.9750 0.3000 ;
        RECT 0.9150 0.8250 0.9750 0.8850 ;
        RECT 0.8100 0.4950 0.8700 0.5550 ;
        RECT 0.7050 0.3075 0.7650 0.3675 ;
        RECT 0.6000 0.4875 0.6600 0.5475 ;
        RECT 0.4950 0.1575 0.5550 0.2175 ;
        RECT 0.4950 0.8025 0.5550 0.8625 ;
        RECT 0.3900 0.4875 0.4500 0.5475 ;
        RECT 0.2850 0.3075 0.3450 0.3675 ;
        RECT 0.1800 0.4950 0.2400 0.5550 ;
        RECT 0.0750 0.1725 0.1350 0.2325 ;
        RECT 0.0750 0.8325 0.1350 0.8925 ;
        LAYER M1 ;
        RECT 2.0700 0.4425 2.7900 0.5475 ;
        RECT 2.5725 0.1950 2.6775 0.3675 ;
        RECT 2.5875 0.6225 2.6625 0.8700 ;
        RECT 2.2425 0.6225 2.5875 0.7125 ;
        RECT 2.2575 0.2775 2.5725 0.3675 ;
        RECT 2.1525 0.1950 2.2575 0.3675 ;
        RECT 2.1675 0.6225 2.2425 0.8700 ;
        RECT 1.9950 0.4425 2.0700 0.6750 ;
        RECT 1.8150 0.4650 1.9200 0.7275 ;
        RECT 0.9900 0.3150 1.8450 0.3900 ;
        RECT 1.3125 0.6525 1.8150 0.7275 ;
        RECT 1.4025 0.8025 1.7475 0.9000 ;
        RECT 1.4100 0.4725 1.7325 0.5775 ;
        RECT 1.2375 0.4725 1.3125 0.7275 ;
        RECT 1.1175 0.4725 1.2375 0.6600 ;
        RECT 0.9150 0.1500 0.9900 0.3900 ;
        RECT 0.1575 0.1500 0.9150 0.2250 ;
        RECT 0.4650 0.7800 0.8400 0.8850 ;
        RECT 0.2475 0.3000 0.8100 0.3750 ;
        RECT 0.3600 0.4500 0.6900 0.5550 ;
        RECT 0.0525 0.1500 0.1575 0.2550 ;
        LAYER VIA1 ;
        RECT 1.9950 0.5475 2.0700 0.6225 ;
        RECT 1.5375 0.8100 1.6125 0.8850 ;
        RECT 0.7275 0.7950 0.8025 0.8700 ;
        RECT 0.6900 0.3000 0.7650 0.3750 ;
        LAYER M2 ;
        RECT 1.9800 0.5100 2.0850 0.8850 ;
        RECT 0.7800 0.7800 1.9800 0.8850 ;
        RECT 0.6750 0.2625 0.7800 0.8850 ;
    END
END OA22_0111


MACRO OA22_1000
    CLASS CORE ;
    FOREIGN OA22_1000 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.4700 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 1.3575 0.1500 1.4325 0.9000 ;
        RECT 1.3125 0.1500 1.3575 0.3825 ;
        RECT 1.3275 0.6675 1.3575 0.9000 ;
        END
    END Z
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.8775 0.4125 1.3425 0.4875 ;
        VIA 0.9900 0.4500 VIA12_square ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.7575 0.1125 1.2075 0.1875 ;
        RECT 0.6525 0.1125 0.7575 0.5700 ;
        VIA 0.7050 0.4875 VIA12_square ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1425 0.5100 0.2700 0.6150 ;
        RECT 0.0675 0.3675 0.1425 0.6825 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.5775 0.7125 1.0950 0.7875 ;
        RECT 0.5025 0.5550 0.5775 0.7875 ;
        VIA 0.5400 0.6750 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.2150 -0.0750 1.4700 0.0750 ;
        RECT 1.0950 -0.0750 1.2150 0.2475 ;
        RECT 0.7950 -0.0750 1.0950 0.0750 ;
        RECT 0.6750 -0.0750 0.7950 0.1800 ;
        RECT 0.0000 -0.0750 0.6750 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.2150 0.9750 1.4700 1.1250 ;
        RECT 1.0950 0.8325 1.2150 1.1250 ;
        RECT 1.0050 0.9750 1.0950 1.1250 ;
        RECT 0.8850 0.8325 1.0050 1.1250 ;
        RECT 0.1650 0.9750 0.8850 1.1250 ;
        RECT 0.0450 0.8025 0.1650 1.1250 ;
        RECT 0.0000 0.9750 0.0450 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.3350 0.1725 1.3950 0.2325 ;
        RECT 1.3350 0.8100 1.3950 0.8700 ;
        RECT 1.2225 0.4950 1.2825 0.5550 ;
        RECT 1.1250 0.1575 1.1850 0.2175 ;
        RECT 1.1250 0.8325 1.1850 0.8925 ;
        RECT 0.9150 0.1725 0.9750 0.2325 ;
        RECT 0.9150 0.8325 0.9750 0.8925 ;
        RECT 0.8175 0.4950 0.8775 0.5550 ;
        RECT 0.7050 0.1200 0.7650 0.1800 ;
        RECT 0.6000 0.4950 0.6600 0.5550 ;
        RECT 0.4950 0.1575 0.5550 0.2175 ;
        RECT 0.4950 0.7950 0.5550 0.8550 ;
        RECT 0.3825 0.5400 0.4425 0.6000 ;
        RECT 0.1800 0.5100 0.2400 0.5700 ;
        RECT 0.0750 0.1650 0.1350 0.2250 ;
        RECT 0.0750 0.8325 0.1350 0.8925 ;
        RECT 0.2850 0.3375 0.3450 0.3975 ;
        LAYER M1 ;
        RECT 1.2525 0.4650 1.2825 0.5850 ;
        RECT 1.1775 0.4650 1.2525 0.7575 ;
        RECT 0.8100 0.6825 1.1775 0.7575 ;
        RECT 0.8175 0.4125 1.0875 0.6000 ;
        RECT 0.8850 0.1500 0.9975 0.3300 ;
        RECT 0.6000 0.2550 0.8850 0.3300 ;
        RECT 0.7350 0.6825 0.8100 0.8625 ;
        RECT 0.6675 0.4050 0.7425 0.5775 ;
        RECT 0.3075 0.7875 0.7350 0.8625 ;
        RECT 0.5475 0.4050 0.6675 0.5625 ;
        RECT 0.4725 0.6375 0.6225 0.7125 ;
        RECT 0.5250 0.1500 0.6000 0.3300 ;
        RECT 0.1500 0.1500 0.5250 0.2250 ;
        RECT 0.3525 0.5400 0.4725 0.7125 ;
        RECT 0.3450 0.3000 0.4500 0.4650 ;
        RECT 0.2175 0.3000 0.3450 0.4350 ;
        RECT 0.0450 0.1500 0.1500 0.2550 ;
        LAYER VIA1 ;
        RECT 0.3525 0.3450 0.4275 0.4200 ;
        RECT 0.3525 0.7875 0.4275 0.8625 ;
        LAYER M2 ;
        RECT 0.4275 0.8625 0.4575 0.9375 ;
        RECT 0.3525 0.3000 0.4275 0.9375 ;
    END
END OA22_1000


MACRO OA22_1010
    CLASS CORE ;
    FOREIGN OA22_1010 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.4700 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 1.3575 0.2175 1.4325 0.8325 ;
        RECT 1.3275 0.2175 1.3575 0.3825 ;
        RECT 1.3275 0.6675 1.3575 0.8325 ;
        END
    END Z
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.8775 0.4125 1.3425 0.4875 ;
        VIA 0.9900 0.4500 VIA12_square ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.7575 0.1125 1.2075 0.1875 ;
        RECT 0.6525 0.1125 0.7575 0.5700 ;
        VIA 0.7050 0.4875 VIA12_square ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1425 0.5100 0.2700 0.6150 ;
        RECT 0.0675 0.3675 0.1425 0.6825 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.5775 0.7125 1.0950 0.7875 ;
        RECT 0.5025 0.5550 0.5775 0.7875 ;
        VIA 0.5400 0.6750 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.2150 -0.0750 1.4700 0.0750 ;
        RECT 1.0950 -0.0750 1.2150 0.2475 ;
        RECT 0.7950 -0.0750 1.0950 0.0750 ;
        RECT 0.6750 -0.0750 0.7950 0.1800 ;
        RECT 0.0000 -0.0750 0.6750 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.2150 0.9750 1.4700 1.1250 ;
        RECT 1.0950 0.8325 1.2150 1.1250 ;
        RECT 1.0050 0.9750 1.0950 1.1250 ;
        RECT 0.8850 0.8325 1.0050 1.1250 ;
        RECT 0.1650 0.9750 0.8850 1.1250 ;
        RECT 0.0450 0.8025 0.1650 1.1250 ;
        RECT 0.0000 0.9750 0.0450 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.3350 0.2700 1.3950 0.3300 ;
        RECT 1.3350 0.7200 1.3950 0.7800 ;
        RECT 1.2225 0.4950 1.2825 0.5550 ;
        RECT 1.1250 0.1575 1.1850 0.2175 ;
        RECT 1.1250 0.8325 1.1850 0.8925 ;
        RECT 0.9150 0.2325 0.9750 0.2925 ;
        RECT 0.9150 0.8325 0.9750 0.8925 ;
        RECT 0.8175 0.4950 0.8775 0.5550 ;
        RECT 0.7050 0.1200 0.7650 0.1800 ;
        RECT 0.6000 0.4950 0.6600 0.5550 ;
        RECT 0.4950 0.1575 0.5550 0.2175 ;
        RECT 0.4950 0.7950 0.5550 0.8550 ;
        RECT 0.3825 0.5400 0.4425 0.6000 ;
        RECT 0.1800 0.5100 0.2400 0.5700 ;
        RECT 0.0750 0.1650 0.1350 0.2250 ;
        RECT 0.0750 0.8325 0.1350 0.8925 ;
        RECT 0.2850 0.3375 0.3450 0.3975 ;
        LAYER M1 ;
        RECT 1.2525 0.4650 1.2825 0.5850 ;
        RECT 1.1775 0.4650 1.2525 0.7575 ;
        RECT 0.8100 0.6825 1.1775 0.7575 ;
        RECT 0.8175 0.4125 1.0875 0.6000 ;
        RECT 0.8850 0.1950 0.9750 0.3300 ;
        RECT 0.6000 0.2550 0.8850 0.3300 ;
        RECT 0.7350 0.6825 0.8100 0.8625 ;
        RECT 0.6675 0.4050 0.7425 0.5775 ;
        RECT 0.3075 0.7875 0.7350 0.8625 ;
        RECT 0.5475 0.4050 0.6675 0.5625 ;
        RECT 0.4725 0.6375 0.6225 0.7125 ;
        RECT 0.5250 0.1500 0.6000 0.3300 ;
        RECT 0.1500 0.1500 0.5250 0.2250 ;
        RECT 0.3525 0.5400 0.4725 0.7125 ;
        RECT 0.3450 0.3000 0.4500 0.4650 ;
        RECT 0.2175 0.3000 0.3450 0.4350 ;
        RECT 0.0450 0.1500 0.1500 0.2550 ;
        LAYER VIA1 ;
        RECT 0.3525 0.3450 0.4275 0.4200 ;
        RECT 0.3525 0.7875 0.4275 0.8625 ;
        LAYER M2 ;
        RECT 0.4275 0.8625 0.4575 0.9375 ;
        RECT 0.3525 0.3000 0.4275 0.9375 ;
    END
END OA22_1010


MACRO OA31_0011
    CLASS CORE ;
    FOREIGN OA31_0011 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.4700 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 1.3575 0.3075 1.4325 0.7425 ;
        RECT 1.1925 0.3075 1.3575 0.3825 ;
        RECT 1.1925 0.6675 1.3575 0.7425 ;
        RECT 1.1175 0.2175 1.1925 0.3825 ;
        RECT 1.1175 0.6675 1.1925 0.8550 ;
        END
    END Z
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.8475 0.8625 1.1925 0.9375 ;
        RECT 0.7725 0.5250 0.8475 0.9375 ;
        RECT 0.6525 0.8625 0.7725 0.9375 ;
        VIA 0.8100 0.6075 VIA12_square ;
        END
    END B
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.6525 0.2625 1.0875 0.3375 ;
        RECT 0.5775 0.2625 0.6525 0.6525 ;
        VIA 0.6150 0.5325 VIA12_square ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.4725 0.1125 0.9225 0.1875 ;
        RECT 0.3675 0.1125 0.4725 0.6150 ;
        VIA 0.4200 0.5325 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.0675 0.7125 0.5325 0.7875 ;
        VIA 0.2550 0.7500 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.4250 -0.0750 1.4700 0.0750 ;
        RECT 1.3050 -0.0750 1.4250 0.2175 ;
        RECT 1.0050 -0.0750 1.3050 0.0750 ;
        RECT 0.9000 -0.0750 1.0050 0.2100 ;
        RECT 0.0000 -0.0750 0.9000 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.4250 0.9750 1.4700 1.1250 ;
        RECT 1.3050 0.8175 1.4250 1.1250 ;
        RECT 1.0050 0.9750 1.3050 1.1250 ;
        RECT 0.8850 0.8700 1.0050 1.1250 ;
        RECT 0.1425 0.9750 0.8850 1.1250 ;
        RECT 0.0675 0.7200 0.1425 1.1250 ;
        RECT 0.0000 0.9750 0.0675 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.3350 0.1575 1.3950 0.2175 ;
        RECT 1.3350 0.8325 1.3950 0.8925 ;
        RECT 1.2225 0.4950 1.2825 0.5550 ;
        RECT 1.1250 0.2775 1.1850 0.3375 ;
        RECT 1.1250 0.7650 1.1850 0.8250 ;
        RECT 1.0200 0.4950 1.0800 0.5550 ;
        RECT 0.9150 0.1200 0.9750 0.1800 ;
        RECT 0.9150 0.8700 0.9750 0.9300 ;
        RECT 0.8100 0.4950 0.8700 0.5550 ;
        RECT 0.7050 0.1575 0.7650 0.2175 ;
        RECT 0.7050 0.7500 0.7650 0.8100 ;
        RECT 0.5925 0.4950 0.6525 0.5550 ;
        RECT 0.4950 0.3075 0.5550 0.3675 ;
        RECT 0.3900 0.4950 0.4500 0.5550 ;
        RECT 0.2850 0.1575 0.3450 0.2175 ;
        RECT 0.1800 0.4950 0.2400 0.5550 ;
        RECT 0.0750 0.2325 0.1350 0.2925 ;
        RECT 0.0750 0.7575 0.1350 0.8175 ;
        LAYER M1 ;
        RECT 1.0425 0.4650 1.2825 0.5850 ;
        RECT 0.9675 0.3000 1.0425 0.7950 ;
        RECT 0.1425 0.3000 0.9675 0.3750 ;
        RECT 0.7725 0.7200 0.9675 0.7950 ;
        RECT 0.7275 0.4500 0.8925 0.6450 ;
        RECT 0.2550 0.1500 0.7950 0.2250 ;
        RECT 0.6975 0.7200 0.7725 0.8400 ;
        RECT 0.6225 0.4500 0.6525 0.6225 ;
        RECT 0.5475 0.4500 0.6225 0.8325 ;
        RECT 0.3675 0.4500 0.4725 0.8325 ;
        RECT 0.2175 0.4500 0.2925 0.8325 ;
        RECT 0.1500 0.4500 0.2175 0.6000 ;
        RECT 0.0675 0.2025 0.1425 0.3750 ;
    END
END OA31_0011


MACRO OA31_0111
    CLASS CORE ;
    FOREIGN OA31_0111 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.7300 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 1.8375 0.2775 2.1525 0.7425 ;
        VIA 1.9950 0.3375 VIA12_slot ;
        VIA 1.9950 0.6825 VIA12_slot ;
        END
    END Z
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 2.3775 0.5625 2.6325 0.6375 ;
        RECT 2.3025 0.5625 2.3775 0.9375 ;
        RECT 1.5300 0.8625 2.3025 0.9375 ;
        RECT 1.4550 0.5625 1.5300 0.9375 ;
        RECT 1.3275 0.5625 1.4550 0.6375 ;
        VIA 2.5500 0.6000 VIA12_square ;
        VIA 1.4400 0.6000 VIA12_square ;
        END
    END B
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.1425 0.7125 1.3050 0.7875 ;
        VIA 1.1925 0.7500 VIA12_square ;
        VIA 0.2550 0.7500 VIA12_square ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.1200 0.5625 0.5850 0.6375 ;
        VIA 0.4575 0.6000 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.8100 0.5625 1.2075 0.6375 ;
        RECT 0.7050 0.4500 0.8100 0.6375 ;
        VIA 0.7575 0.5250 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 2.4750 -0.0750 2.7300 0.0750 ;
        RECT 2.3550 -0.0750 2.4750 0.1800 ;
        RECT 2.0550 -0.0750 2.3550 0.0750 ;
        RECT 1.9350 -0.0750 2.0550 0.1950 ;
        RECT 1.6350 -0.0750 1.9350 0.0750 ;
        RECT 1.5150 -0.0750 1.6350 0.1875 ;
        RECT 0.0000 -0.0750 1.5150 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 2.4750 0.9750 2.7300 1.1250 ;
        RECT 2.3550 0.8700 2.4750 1.1250 ;
        RECT 2.0550 0.9750 2.3550 1.1250 ;
        RECT 1.9350 0.8625 2.0550 1.1250 ;
        RECT 1.6350 0.9750 1.9350 1.1250 ;
        RECT 1.5150 0.8700 1.6350 1.1250 ;
        RECT 0.7950 0.9750 1.5150 1.1250 ;
        RECT 0.6750 0.8250 0.7950 1.1250 ;
        RECT 0.0000 0.9750 0.6750 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 2.5950 0.2250 2.6550 0.2850 ;
        RECT 2.5950 0.7500 2.6550 0.8100 ;
        RECT 2.4900 0.4950 2.5500 0.5550 ;
        RECT 2.3850 0.1200 2.4450 0.1800 ;
        RECT 2.3850 0.8700 2.4450 0.9300 ;
        RECT 2.2800 0.4650 2.3400 0.5250 ;
        RECT 2.1750 0.2250 2.2350 0.2850 ;
        RECT 2.1750 0.7575 2.2350 0.8175 ;
        RECT 2.0700 0.4650 2.1300 0.5250 ;
        RECT 1.9650 0.1275 2.0250 0.1875 ;
        RECT 1.9650 0.8700 2.0250 0.9300 ;
        RECT 1.8600 0.4650 1.9200 0.5250 ;
        RECT 1.7550 0.2250 1.8150 0.2850 ;
        RECT 1.7550 0.7575 1.8150 0.8175 ;
        RECT 1.6500 0.4650 1.7100 0.5250 ;
        RECT 1.5450 0.1275 1.6050 0.1875 ;
        RECT 1.5450 0.8700 1.6050 0.9300 ;
        RECT 1.4400 0.4950 1.5000 0.5550 ;
        RECT 1.3350 0.1575 1.3950 0.2175 ;
        RECT 1.3350 0.7575 1.3950 0.8175 ;
        RECT 1.2225 0.4950 1.2825 0.5550 ;
        RECT 1.1250 0.3075 1.1850 0.3675 ;
        RECT 1.0200 0.4950 1.0800 0.5550 ;
        RECT 0.9150 0.1575 0.9750 0.2175 ;
        RECT 0.8100 0.4875 0.8700 0.5475 ;
        RECT 0.7050 0.3075 0.7650 0.3675 ;
        RECT 0.7050 0.8475 0.7650 0.9075 ;
        RECT 0.6000 0.4875 0.6600 0.5475 ;
        RECT 0.4950 0.1575 0.5550 0.2175 ;
        RECT 0.3900 0.4950 0.4500 0.5550 ;
        RECT 0.2850 0.3075 0.3450 0.3675 ;
        RECT 0.1875 0.5100 0.2475 0.5700 ;
        RECT 0.0750 0.1725 0.1350 0.2325 ;
        RECT 0.0750 0.7800 0.1350 0.8400 ;
        LAYER M1 ;
        RECT 2.5875 0.1875 2.6625 0.3600 ;
        RECT 2.4675 0.4350 2.6625 0.6450 ;
        RECT 2.5875 0.7200 2.6625 0.8400 ;
        RECT 2.3175 0.2550 2.5875 0.3600 ;
        RECT 2.3925 0.7200 2.5875 0.7950 ;
        RECT 2.3175 0.4575 2.3925 0.7950 ;
        RECT 1.6725 0.4575 2.3175 0.5475 ;
        RECT 2.1675 0.1950 2.2425 0.3825 ;
        RECT 2.1675 0.6225 2.2425 0.8700 ;
        RECT 1.8375 0.2925 2.1675 0.3825 ;
        RECT 1.8225 0.6225 2.1675 0.7425 ;
        RECT 1.7325 0.1950 1.8375 0.3825 ;
        RECT 1.7475 0.6225 1.8225 0.8700 ;
        RECT 1.5975 0.4575 1.6725 0.7950 ;
        RECT 1.4025 0.7200 1.5975 0.7950 ;
        RECT 1.4400 0.2625 1.5900 0.3375 ;
        RECT 1.3575 0.4500 1.5225 0.6450 ;
        RECT 1.3500 0.1500 1.4400 0.3375 ;
        RECT 1.3275 0.7200 1.4025 0.8550 ;
        RECT 0.1575 0.1500 1.3500 0.2250 ;
        RECT 1.2300 0.4500 1.2825 0.5850 ;
        RECT 0.3300 0.3000 1.2375 0.3750 ;
        RECT 1.1550 0.4500 1.2300 0.8475 ;
        RECT 0.9750 0.4650 1.0800 0.7200 ;
        RECT 0.4950 0.6450 0.9750 0.7200 ;
        RECT 0.5700 0.4650 0.9000 0.5700 ;
        RECT 0.4200 0.4650 0.4950 0.7200 ;
        RECT 0.3825 0.4650 0.4200 0.5850 ;
        RECT 0.2925 0.7950 0.3900 0.9000 ;
        RECT 0.2550 0.3000 0.3300 0.4050 ;
        RECT 0.2100 0.4800 0.2925 0.9000 ;
        RECT 0.1125 0.3300 0.2550 0.4050 ;
        RECT 0.1875 0.4800 0.2100 0.6600 ;
        RECT 0.0525 0.1500 0.1575 0.2550 ;
        RECT 0.1125 0.7500 0.1350 0.8700 ;
        RECT 0.0375 0.3300 0.1125 0.8700 ;
        LAYER VIA1 ;
        RECT 2.3625 0.2625 2.4375 0.3375 ;
        RECT 1.6425 0.4650 1.7175 0.5400 ;
        RECT 1.4400 0.2625 1.5150 0.3375 ;
        RECT 1.0800 0.3000 1.1550 0.3750 ;
        LAYER M2 ;
        RECT 2.3625 0.2625 2.4825 0.3375 ;
        RECT 2.2800 0.1125 2.3625 0.3375 ;
        RECT 1.7025 0.1125 2.2800 0.1875 ;
        RECT 1.6275 0.4125 1.7325 0.5775 ;
        RECT 1.6275 0.1125 1.7025 0.3375 ;
        RECT 1.3650 0.2625 1.6275 0.3375 ;
        RECT 1.2450 0.4125 1.6275 0.4875 ;
        RECT 1.1700 0.3000 1.2450 0.4875 ;
        RECT 1.0050 0.3000 1.1700 0.3750 ;
    END
END OA31_0111


MACRO OA31_1000
    CLASS CORE ;
    FOREIGN OA31_1000 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.2600 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 1.1475 0.1500 1.2225 0.9000 ;
        RECT 1.1175 0.1500 1.1475 0.3825 ;
        RECT 1.1175 0.6675 1.1475 0.9000 ;
        END
    END Z
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.8475 0.8625 1.1925 0.9375 ;
        RECT 0.7725 0.5250 0.8475 0.9375 ;
        RECT 0.6525 0.8625 0.7725 0.9375 ;
        VIA 0.8100 0.6075 VIA12_square ;
        END
    END B
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.6525 0.2625 1.0875 0.3375 ;
        RECT 0.5775 0.2625 0.6525 0.6525 ;
        VIA 0.6150 0.5325 VIA12_square ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.4725 0.1125 0.9225 0.1875 ;
        RECT 0.3675 0.1125 0.4725 0.6150 ;
        VIA 0.4200 0.5325 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.0675 0.7125 0.5325 0.7875 ;
        VIA 0.2550 0.7500 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.0050 -0.0750 1.2600 0.0750 ;
        RECT 0.9000 -0.0750 1.0050 0.2100 ;
        RECT 0.0000 -0.0750 0.9000 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.0050 0.9750 1.2600 1.1250 ;
        RECT 0.8850 0.8700 1.0050 1.1250 ;
        RECT 0.1425 0.9750 0.8850 1.1250 ;
        RECT 0.0675 0.7950 0.1425 1.1250 ;
        RECT 0.0000 0.9750 0.0675 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.1250 0.1800 1.1850 0.2400 ;
        RECT 1.1250 0.8100 1.1850 0.8700 ;
        RECT 1.0125 0.4950 1.0725 0.5550 ;
        RECT 0.9150 0.1200 0.9750 0.1800 ;
        RECT 0.9150 0.8700 0.9750 0.9300 ;
        RECT 0.8100 0.4950 0.8700 0.5550 ;
        RECT 0.7050 0.1575 0.7650 0.2175 ;
        RECT 0.7050 0.7800 0.7650 0.8400 ;
        RECT 0.5925 0.4950 0.6525 0.5550 ;
        RECT 0.4950 0.3000 0.5550 0.3600 ;
        RECT 0.3900 0.4950 0.4500 0.5550 ;
        RECT 0.2850 0.1575 0.3450 0.2175 ;
        RECT 0.1800 0.4950 0.2400 0.5550 ;
        RECT 0.0750 0.2325 0.1350 0.2925 ;
        RECT 0.0750 0.8325 0.1350 0.8925 ;
        LAYER M1 ;
        RECT 1.0425 0.4650 1.0725 0.5850 ;
        RECT 0.9675 0.3000 1.0425 0.7950 ;
        RECT 0.1425 0.3000 0.9675 0.3750 ;
        RECT 0.7725 0.7200 0.9675 0.7950 ;
        RECT 0.7275 0.4500 0.8925 0.6450 ;
        RECT 0.2550 0.1500 0.7950 0.2250 ;
        RECT 0.6975 0.7200 0.7725 0.8700 ;
        RECT 0.6225 0.4500 0.6525 0.6225 ;
        RECT 0.5475 0.4500 0.6225 0.8325 ;
        RECT 0.3675 0.4500 0.4725 0.8325 ;
        RECT 0.2175 0.4500 0.2925 0.8325 ;
        RECT 0.1500 0.4500 0.2175 0.6000 ;
        RECT 0.0675 0.2025 0.1425 0.3750 ;
    END
END OA31_1000


MACRO OA31_1010
    CLASS CORE ;
    FOREIGN OA31_1010 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.2600 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 1.1475 0.2175 1.2225 0.8325 ;
        RECT 1.1175 0.2175 1.1475 0.3825 ;
        RECT 1.1175 0.6675 1.1475 0.8325 ;
        END
    END Z
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.8475 0.8625 1.1925 0.9375 ;
        RECT 0.7725 0.5250 0.8475 0.9375 ;
        RECT 0.6525 0.8625 0.7725 0.9375 ;
        VIA 0.8100 0.6075 VIA12_square ;
        END
    END B
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.6525 0.2625 1.0875 0.3375 ;
        RECT 0.5775 0.2625 0.6525 0.6525 ;
        VIA 0.6150 0.5325 VIA12_square ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.4725 0.1125 0.9225 0.1875 ;
        RECT 0.3675 0.1125 0.4725 0.6150 ;
        VIA 0.4200 0.5325 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.0675 0.7125 0.5325 0.7875 ;
        VIA 0.2550 0.7500 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.0050 -0.0750 1.2600 0.0750 ;
        RECT 0.9000 -0.0750 1.0050 0.2100 ;
        RECT 0.0000 -0.0750 0.9000 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.0050 0.9750 1.2600 1.1250 ;
        RECT 0.8850 0.8700 1.0050 1.1250 ;
        RECT 0.1425 0.9750 0.8850 1.1250 ;
        RECT 0.0675 0.7200 0.1425 1.1250 ;
        RECT 0.0000 0.9750 0.0675 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.1250 0.2625 1.1850 0.3225 ;
        RECT 1.1250 0.7200 1.1850 0.7800 ;
        RECT 1.0125 0.4950 1.0725 0.5550 ;
        RECT 0.9150 0.1200 0.9750 0.1800 ;
        RECT 0.9150 0.8700 0.9750 0.9300 ;
        RECT 0.8100 0.4950 0.8700 0.5550 ;
        RECT 0.7050 0.1575 0.7650 0.2175 ;
        RECT 0.7050 0.7500 0.7650 0.8100 ;
        RECT 0.5925 0.4950 0.6525 0.5550 ;
        RECT 0.4950 0.3075 0.5550 0.3675 ;
        RECT 0.3900 0.4950 0.4500 0.5550 ;
        RECT 0.2850 0.1575 0.3450 0.2175 ;
        RECT 0.1800 0.4950 0.2400 0.5550 ;
        RECT 0.0750 0.2325 0.1350 0.2925 ;
        RECT 0.0750 0.7575 0.1350 0.8175 ;
        LAYER M1 ;
        RECT 1.0425 0.4650 1.0725 0.5850 ;
        RECT 0.9675 0.3000 1.0425 0.7950 ;
        RECT 0.1425 0.3000 0.9675 0.3750 ;
        RECT 0.7725 0.7200 0.9675 0.7950 ;
        RECT 0.7275 0.4500 0.8925 0.6450 ;
        RECT 0.2550 0.1500 0.7950 0.2250 ;
        RECT 0.6975 0.7200 0.7725 0.8400 ;
        RECT 0.6225 0.4500 0.6525 0.6225 ;
        RECT 0.5475 0.4500 0.6225 0.8325 ;
        RECT 0.3675 0.4500 0.4725 0.8325 ;
        RECT 0.2175 0.4500 0.2925 0.8325 ;
        RECT 0.1500 0.4500 0.2175 0.6000 ;
        RECT 0.0675 0.2025 0.1425 0.3750 ;
    END
END OA31_1010


MACRO OA32_0011
    CLASS CORE ;
    FOREIGN OA32_0011 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.8900 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.2775 0.2175 0.3525 0.3675 ;
        RECT 0.2775 0.6675 0.3525 0.8550 ;
        RECT 0.1125 0.2925 0.2775 0.3675 ;
        RECT 0.1125 0.6675 0.2775 0.7425 ;
        RECT 0.0375 0.2925 0.1125 0.7425 ;
        END
    END Z
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.3575 0.7125 1.8225 0.7875 ;
        VIA 1.5150 0.7500 VIA12_square ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.3575 0.5625 1.8225 0.6375 ;
        VIA 1.6800 0.6000 VIA12_square ;
        END
    END B1
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.2375 0.1125 1.8225 0.1875 ;
        RECT 1.1625 0.1125 1.2375 0.6600 ;
        VIA 1.2000 0.5325 VIA12_square ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.9675 0.1125 1.0425 0.6600 ;
        RECT 0.5175 0.1125 0.9675 0.1875 ;
        RECT 0.9150 0.5550 0.9675 0.6600 ;
        VIA 1.0050 0.5175 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.7425 0.4575 0.8175 0.6375 ;
        RECT 0.2775 0.5625 0.7425 0.6375 ;
        VIA 0.7800 0.5400 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.6350 -0.0750 1.8900 0.0750 ;
        RECT 1.5150 -0.0750 1.6350 0.1950 ;
        RECT 0.5850 -0.0750 1.5150 0.0750 ;
        RECT 0.4650 -0.0750 0.5850 0.2250 ;
        RECT 0.1650 -0.0750 0.4650 0.0750 ;
        RECT 0.0450 -0.0750 0.1650 0.2175 ;
        RECT 0.0000 -0.0750 0.0450 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.8450 0.9750 1.8900 1.1250 ;
        RECT 1.7250 0.7875 1.8450 1.1250 ;
        RECT 0.7875 0.9750 1.7250 1.1250 ;
        RECT 0.6825 0.8100 0.7875 1.1250 ;
        RECT 0.5775 0.9750 0.6825 1.1250 ;
        RECT 0.4725 0.8100 0.5775 1.1250 ;
        RECT 0.1650 0.9750 0.4725 1.1250 ;
        RECT 0.0450 0.8175 0.1650 1.1250 ;
        RECT 0.0000 0.9750 0.0450 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.7550 0.2475 1.8150 0.3075 ;
        RECT 1.7550 0.8175 1.8150 0.8775 ;
        RECT 1.6500 0.4950 1.7100 0.5550 ;
        RECT 1.5450 0.1350 1.6050 0.1950 ;
        RECT 1.4400 0.4950 1.5000 0.5550 ;
        RECT 1.3350 0.1575 1.3950 0.2175 ;
        RECT 1.3350 0.8100 1.3950 0.8700 ;
        RECT 1.2300 0.4950 1.2900 0.5550 ;
        RECT 1.1250 0.3075 1.1850 0.3675 ;
        RECT 1.0200 0.4950 1.0800 0.5550 ;
        RECT 0.9150 0.1575 0.9750 0.2175 ;
        RECT 0.8025 0.4875 0.8625 0.5475 ;
        RECT 0.7050 0.3000 0.7650 0.3600 ;
        RECT 0.7050 0.8325 0.7650 0.8925 ;
        RECT 0.4950 0.1575 0.5550 0.2175 ;
        RECT 0.4950 0.8325 0.5550 0.8925 ;
        RECT 0.3900 0.4950 0.4500 0.5550 ;
        RECT 0.2850 0.2550 0.3450 0.3150 ;
        RECT 0.2850 0.7650 0.3450 0.8250 ;
        RECT 0.1875 0.4950 0.2475 0.5550 ;
        RECT 0.0750 0.1575 0.1350 0.2175 ;
        RECT 0.0750 0.8325 0.1350 0.8925 ;
        LAYER M1 ;
        RECT 1.7400 0.2175 1.8300 0.3450 ;
        RECT 1.6425 0.4575 1.7925 0.6825 ;
        RECT 1.4400 0.2700 1.7400 0.3450 ;
        RECT 1.6200 0.4575 1.6425 0.5625 ;
        RECT 1.5450 0.6450 1.5675 0.8325 ;
        RECT 1.4700 0.4200 1.5450 0.8325 ;
        RECT 1.4400 0.4200 1.4700 0.7200 ;
        RECT 1.3650 0.1500 1.4400 0.3450 ;
        RECT 1.2900 0.7800 1.3950 0.9000 ;
        RECT 0.8850 0.1500 1.3650 0.2250 ;
        RECT 1.1625 0.4500 1.3650 0.6150 ;
        RECT 0.9375 0.8250 1.2900 0.9000 ;
        RECT 0.5025 0.3000 1.2150 0.3750 ;
        RECT 1.0875 0.6750 1.1175 0.7500 ;
        RECT 1.0125 0.4500 1.0875 0.7500 ;
        RECT 0.9375 0.4500 1.0125 0.5850 ;
        RECT 0.8625 0.6600 0.9375 0.9000 ;
        RECT 0.5775 0.4500 0.8625 0.5775 ;
        RECT 0.5025 0.6600 0.8625 0.7350 ;
        RECT 0.4275 0.3000 0.5025 0.7350 ;
        RECT 0.1875 0.4650 0.4275 0.5850 ;
    END
END OA32_0011


MACRO OA32_0111
    CLASS CORE ;
    FOREIGN OA32_0111 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.3600 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 2.6775 0.2400 2.9925 0.7500 ;
        VIA 2.8350 0.3225 VIA12_slot ;
        VIA 2.8350 0.6675 VIA12_slot ;
        END
    END Z
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.5175 0.4425 0.6225 0.7875 ;
        RECT 0.0975 0.7125 0.5175 0.7875 ;
        VIA 0.5700 0.5250 VIA12_square ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.7650 0.2625 0.8700 0.5775 ;
        RECT 0.4275 0.2625 0.7650 0.3375 ;
        RECT 0.3525 0.2625 0.4275 0.4875 ;
        RECT 0.1425 0.4125 0.3525 0.4875 ;
        VIA 0.8175 0.4950 VIA12_square ;
        VIA 0.2250 0.4500 VIA12_square ;
        END
    END B1
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.5375 0.2625 1.6425 0.6225 ;
        RECT 1.0650 0.2625 1.5375 0.3375 ;
        VIA 1.5900 0.5250 VIA12_square ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.8075 0.1125 1.9125 0.6300 ;
        RECT 1.3350 0.1125 1.8075 0.1875 ;
        VIA 1.8600 0.5475 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 2.0325 0.4425 2.1225 0.7875 ;
        RECT 1.1625 0.7125 2.0325 0.7875 ;
        RECT 1.0575 0.4725 1.1625 0.7875 ;
        VIA 2.0775 0.5250 VIA12_square ;
        VIA 1.1100 0.5550 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 3.2925 -0.0750 3.3600 0.0750 ;
        RECT 3.2175 -0.0750 3.2925 0.3150 ;
        RECT 2.8950 -0.0750 3.2175 0.0750 ;
        RECT 2.7750 -0.0750 2.8950 0.1950 ;
        RECT 2.4750 -0.0750 2.7750 0.0750 ;
        RECT 2.3700 -0.0750 2.4750 0.2475 ;
        RECT 0.7950 -0.0750 2.3700 0.0750 ;
        RECT 0.6750 -0.0750 0.7950 0.1875 ;
        RECT 0.3750 -0.0750 0.6750 0.0750 ;
        RECT 0.2550 -0.0750 0.3750 0.1875 ;
        RECT 0.0000 -0.0750 0.2550 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 3.2925 0.9750 3.3600 1.1250 ;
        RECT 3.2175 0.6375 3.2925 1.1250 ;
        RECT 2.8875 0.9750 3.2175 1.1250 ;
        RECT 2.7825 0.7950 2.8875 1.1250 ;
        RECT 2.4750 0.9750 2.7825 1.1250 ;
        RECT 2.3550 0.8100 2.4750 1.1250 ;
        RECT 2.2650 0.9750 2.3550 1.1250 ;
        RECT 2.1450 0.8100 2.2650 1.1250 ;
        RECT 1.0050 0.9750 2.1450 1.1250 ;
        RECT 0.8850 0.8625 1.0050 1.1250 ;
        RECT 0.1650 0.9750 0.8850 1.1250 ;
        RECT 0.0450 0.6600 0.1650 1.1250 ;
        RECT 0.0000 0.9750 0.0450 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 3.2250 0.2250 3.2850 0.2850 ;
        RECT 3.2250 0.6675 3.2850 0.7275 ;
        RECT 3.2250 0.8325 3.2850 0.8925 ;
        RECT 3.1200 0.4650 3.1800 0.5250 ;
        RECT 3.0150 0.2250 3.0750 0.2850 ;
        RECT 3.0150 0.7575 3.0750 0.8175 ;
        RECT 2.9100 0.4650 2.9700 0.5250 ;
        RECT 2.8050 0.1275 2.8650 0.1875 ;
        RECT 2.8050 0.8250 2.8650 0.8850 ;
        RECT 2.7000 0.4650 2.7600 0.5250 ;
        RECT 2.5950 0.2250 2.6550 0.2850 ;
        RECT 2.5950 0.7575 2.6550 0.8175 ;
        RECT 2.4900 0.4650 2.5500 0.5250 ;
        RECT 2.3850 0.1575 2.4450 0.2175 ;
        RECT 2.3850 0.8175 2.4450 0.8775 ;
        RECT 2.1750 0.1725 2.2350 0.2325 ;
        RECT 2.1750 0.8175 2.2350 0.8775 ;
        RECT 2.0700 0.4950 2.1300 0.5550 ;
        RECT 1.9650 0.3225 2.0250 0.3825 ;
        RECT 1.8600 0.4950 1.9200 0.5550 ;
        RECT 1.7550 0.1725 1.8150 0.2325 ;
        RECT 1.6500 0.4950 1.7100 0.5550 ;
        RECT 1.5450 0.3225 1.6050 0.3825 ;
        RECT 1.5450 0.8175 1.6050 0.8775 ;
        RECT 1.4400 0.4950 1.5000 0.5550 ;
        RECT 1.3350 0.1725 1.3950 0.2325 ;
        RECT 1.2300 0.4950 1.2900 0.5550 ;
        RECT 1.1250 0.3225 1.1850 0.3825 ;
        RECT 1.0200 0.4950 1.0800 0.5550 ;
        RECT 0.9150 0.2250 0.9750 0.2850 ;
        RECT 0.9150 0.8700 0.9750 0.9300 ;
        RECT 0.8100 0.4875 0.8700 0.5475 ;
        RECT 0.7050 0.1200 0.7650 0.1800 ;
        RECT 0.6000 0.4950 0.6600 0.5550 ;
        RECT 0.4950 0.2700 0.5550 0.3300 ;
        RECT 0.4950 0.7200 0.5550 0.7800 ;
        RECT 0.3900 0.4950 0.4500 0.5550 ;
        RECT 0.2850 0.1200 0.3450 0.1800 ;
        RECT 0.1800 0.4725 0.2400 0.5325 ;
        RECT 0.0750 0.2475 0.1350 0.3075 ;
        RECT 0.0750 0.6675 0.1350 0.7275 ;
        RECT 0.0750 0.8325 0.1350 0.8925 ;
        LAYER M1 ;
        RECT 2.4900 0.4425 3.2100 0.5475 ;
        RECT 2.9925 0.1950 3.0975 0.3675 ;
        RECT 3.0075 0.6225 3.0825 0.8700 ;
        RECT 2.6625 0.6225 3.0075 0.7125 ;
        RECT 2.6775 0.2775 2.9925 0.3675 ;
        RECT 2.5725 0.1950 2.6775 0.3675 ;
        RECT 2.5875 0.6225 2.6625 0.8700 ;
        RECT 2.4150 0.3225 2.4900 0.7350 ;
        RECT 2.2800 0.3225 2.4150 0.3975 ;
        RECT 2.0700 0.6600 2.4150 0.7350 ;
        RECT 2.0025 0.4725 2.3025 0.5775 ;
        RECT 2.2125 0.3150 2.2800 0.3975 ;
        RECT 0.9825 0.1650 2.2650 0.2400 ;
        RECT 1.0875 0.3150 2.2125 0.3900 ;
        RECT 1.9950 0.6600 2.0700 0.8850 ;
        RECT 1.1550 0.8100 1.9950 0.8850 ;
        RECT 1.8150 0.4650 1.9200 0.7275 ;
        RECT 1.3350 0.6525 1.8150 0.7275 ;
        RECT 1.4100 0.4725 1.7400 0.5775 ;
        RECT 1.2300 0.4650 1.3350 0.7275 ;
        RECT 0.9600 0.4725 1.1550 0.6375 ;
        RECT 1.0800 0.7125 1.1550 0.8850 ;
        RECT 0.4650 0.7125 1.0800 0.7875 ;
        RECT 0.9075 0.1650 0.9825 0.3375 ;
        RECT 0.1425 0.2625 0.9075 0.3375 ;
        RECT 0.7425 0.4125 0.8850 0.6375 ;
        RECT 0.3825 0.4650 0.6675 0.5850 ;
        RECT 0.1125 0.4125 0.3075 0.5850 ;
        RECT 0.0675 0.2175 0.1425 0.3375 ;
    END
END OA32_0111


MACRO OA32_1000
    CLASS CORE ;
    FOREIGN OA32_1000 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.6800 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1125 0.1500 0.1425 0.3825 ;
        RECT 0.1125 0.6675 0.1425 0.9000 ;
        RECT 0.0375 0.1500 0.1125 0.9000 ;
        END
    END Z
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.1475 0.7125 1.6125 0.7875 ;
        VIA 1.3050 0.7500 VIA12_square ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.1475 0.5625 1.6125 0.6375 ;
        VIA 1.4700 0.6000 VIA12_square ;
        END
    END B1
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.0275 0.1125 1.6125 0.1875 ;
        RECT 0.9525 0.1125 1.0275 0.6600 ;
        VIA 0.9900 0.5325 VIA12_square ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.7575 0.1125 0.8325 0.6600 ;
        RECT 0.3075 0.1125 0.7575 0.1875 ;
        RECT 0.7050 0.5550 0.7575 0.6600 ;
        VIA 0.7950 0.5175 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.5325 0.4575 0.6075 0.6375 ;
        RECT 0.0675 0.5625 0.5325 0.6375 ;
        VIA 0.5700 0.5400 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.4250 -0.0750 1.6800 0.0750 ;
        RECT 1.3050 -0.0750 1.4250 0.1950 ;
        RECT 0.3750 -0.0750 1.3050 0.0750 ;
        RECT 0.2550 -0.0750 0.3750 0.2250 ;
        RECT 0.0000 -0.0750 0.2550 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.6350 0.9750 1.6800 1.1250 ;
        RECT 1.5150 0.7875 1.6350 1.1250 ;
        RECT 0.5775 0.9750 1.5150 1.1250 ;
        RECT 0.4725 0.8100 0.5775 1.1250 ;
        RECT 0.3675 0.9750 0.4725 1.1250 ;
        RECT 0.2625 0.8100 0.3675 1.1250 ;
        RECT 0.0000 0.9750 0.2625 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.5450 0.2475 1.6050 0.3075 ;
        RECT 1.5450 0.8175 1.6050 0.8775 ;
        RECT 1.4400 0.4950 1.5000 0.5550 ;
        RECT 1.3350 0.1350 1.3950 0.1950 ;
        RECT 1.2300 0.4950 1.2900 0.5550 ;
        RECT 1.1250 0.1575 1.1850 0.2175 ;
        RECT 1.1250 0.8100 1.1850 0.8700 ;
        RECT 1.0200 0.4950 1.0800 0.5550 ;
        RECT 0.9150 0.3075 0.9750 0.3675 ;
        RECT 0.8100 0.4950 0.8700 0.5550 ;
        RECT 0.7050 0.1575 0.7650 0.2175 ;
        RECT 0.5925 0.4875 0.6525 0.5475 ;
        RECT 0.4950 0.2250 0.5550 0.2850 ;
        RECT 0.4950 0.8325 0.5550 0.8925 ;
        RECT 0.2850 0.1575 0.3450 0.2175 ;
        RECT 0.2850 0.8325 0.3450 0.8925 ;
        RECT 0.1875 0.4950 0.2475 0.5550 ;
        RECT 0.0750 0.1800 0.1350 0.2400 ;
        RECT 0.0750 0.8100 0.1350 0.8700 ;
        LAYER M1 ;
        RECT 1.5300 0.2175 1.6200 0.3450 ;
        RECT 1.4325 0.4575 1.5825 0.6825 ;
        RECT 1.2300 0.2700 1.5300 0.3450 ;
        RECT 1.4100 0.4575 1.4325 0.5625 ;
        RECT 1.3350 0.6450 1.3575 0.8325 ;
        RECT 1.2600 0.4200 1.3350 0.8325 ;
        RECT 1.2300 0.4200 1.2600 0.7200 ;
        RECT 1.1550 0.1500 1.2300 0.3450 ;
        RECT 1.0800 0.7800 1.1850 0.9000 ;
        RECT 0.6750 0.1500 1.1550 0.2250 ;
        RECT 0.9525 0.4500 1.1550 0.6150 ;
        RECT 0.7275 0.8250 1.0800 0.9000 ;
        RECT 0.5625 0.3000 1.0050 0.3750 ;
        RECT 0.8775 0.6750 0.9075 0.7500 ;
        RECT 0.8025 0.4500 0.8775 0.7500 ;
        RECT 0.7275 0.4500 0.8025 0.5850 ;
        RECT 0.6525 0.6600 0.7275 0.9000 ;
        RECT 0.3675 0.4500 0.6525 0.5775 ;
        RECT 0.2925 0.6600 0.6525 0.7350 ;
        RECT 0.4875 0.1800 0.5625 0.3750 ;
        RECT 0.2925 0.3000 0.4875 0.3750 ;
        RECT 0.2175 0.3000 0.2925 0.7350 ;
        RECT 0.1875 0.4650 0.2175 0.5850 ;
    END
END OA32_1000


MACRO OA32_1010
    CLASS CORE ;
    FOREIGN OA32_1010 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.6800 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1125 0.2175 0.1425 0.3825 ;
        RECT 0.1125 0.6675 0.1425 0.8325 ;
        RECT 0.0375 0.2175 0.1125 0.8325 ;
        END
    END Z
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.1475 0.7125 1.6125 0.7875 ;
        VIA 1.3050 0.7500 VIA12_square ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.1475 0.5625 1.6125 0.6375 ;
        VIA 1.4700 0.6000 VIA12_square ;
        END
    END B1
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.0275 0.1125 1.6125 0.1875 ;
        RECT 0.9525 0.1125 1.0275 0.6600 ;
        VIA 0.9900 0.5325 VIA12_square ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.7575 0.1125 0.8325 0.6600 ;
        RECT 0.3075 0.1125 0.7575 0.1875 ;
        RECT 0.7050 0.5550 0.7575 0.6600 ;
        VIA 0.7950 0.5175 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.5325 0.4575 0.6075 0.6375 ;
        RECT 0.0675 0.5625 0.5325 0.6375 ;
        VIA 0.5700 0.5400 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.4250 -0.0750 1.6800 0.0750 ;
        RECT 1.3050 -0.0750 1.4250 0.1950 ;
        RECT 0.3750 -0.0750 1.3050 0.0750 ;
        RECT 0.2550 -0.0750 0.3750 0.2250 ;
        RECT 0.0000 -0.0750 0.2550 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.6350 0.9750 1.6800 1.1250 ;
        RECT 1.5150 0.7875 1.6350 1.1250 ;
        RECT 0.5775 0.9750 1.5150 1.1250 ;
        RECT 0.4725 0.8100 0.5775 1.1250 ;
        RECT 0.3675 0.9750 0.4725 1.1250 ;
        RECT 0.2625 0.8100 0.3675 1.1250 ;
        RECT 0.0000 0.9750 0.2625 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.5450 0.2475 1.6050 0.3075 ;
        RECT 1.5450 0.8175 1.6050 0.8775 ;
        RECT 1.4400 0.4950 1.5000 0.5550 ;
        RECT 1.3350 0.1350 1.3950 0.1950 ;
        RECT 1.2300 0.4950 1.2900 0.5550 ;
        RECT 1.1250 0.1575 1.1850 0.2175 ;
        RECT 1.1250 0.8100 1.1850 0.8700 ;
        RECT 1.0200 0.4950 1.0800 0.5550 ;
        RECT 0.9150 0.3075 0.9750 0.3675 ;
        RECT 0.8100 0.4950 0.8700 0.5550 ;
        RECT 0.7050 0.1575 0.7650 0.2175 ;
        RECT 0.5925 0.4875 0.6525 0.5475 ;
        RECT 0.4950 0.3000 0.5550 0.3600 ;
        RECT 0.4950 0.8325 0.5550 0.8925 ;
        RECT 0.2850 0.1575 0.3450 0.2175 ;
        RECT 0.2850 0.8325 0.3450 0.8925 ;
        RECT 0.1875 0.4950 0.2475 0.5550 ;
        RECT 0.0750 0.2700 0.1350 0.3300 ;
        RECT 0.0750 0.7200 0.1350 0.7800 ;
        LAYER M1 ;
        RECT 1.5300 0.2175 1.6200 0.3450 ;
        RECT 1.4325 0.4575 1.5825 0.6825 ;
        RECT 1.2300 0.2700 1.5300 0.3450 ;
        RECT 1.4100 0.4575 1.4325 0.5625 ;
        RECT 1.3350 0.6450 1.3575 0.8325 ;
        RECT 1.2600 0.4200 1.3350 0.8325 ;
        RECT 1.2300 0.4200 1.2600 0.7200 ;
        RECT 1.1550 0.1500 1.2300 0.3450 ;
        RECT 1.0800 0.7800 1.1850 0.9000 ;
        RECT 0.6750 0.1500 1.1550 0.2250 ;
        RECT 0.9525 0.4500 1.1550 0.6150 ;
        RECT 0.7275 0.8250 1.0800 0.9000 ;
        RECT 0.2925 0.3000 1.0050 0.3750 ;
        RECT 0.8775 0.6750 0.9075 0.7500 ;
        RECT 0.8025 0.4500 0.8775 0.7500 ;
        RECT 0.7275 0.4500 0.8025 0.5850 ;
        RECT 0.6525 0.6600 0.7275 0.9000 ;
        RECT 0.3675 0.4500 0.6525 0.5775 ;
        RECT 0.2925 0.6600 0.6525 0.7350 ;
        RECT 0.2175 0.3000 0.2925 0.7350 ;
        RECT 0.1875 0.4650 0.2175 0.5850 ;
    END
END OA32_1010


MACRO OA33_0011
    CLASS CORE ;
    FOREIGN OA33_0011 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.8900 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 1.7775 0.3075 1.8525 0.7425 ;
        RECT 1.6125 0.3075 1.7775 0.3825 ;
        RECT 1.6125 0.6675 1.7775 0.7425 ;
        RECT 1.5375 0.2175 1.6125 0.3825 ;
        RECT 1.5375 0.6675 1.6125 0.8550 ;
        END
    END Z
    PIN B3
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.8625 0.4125 1.3200 0.4875 ;
        RECT 0.7575 0.4125 0.8625 0.5850 ;
        VIA 0.8100 0.5025 VIA12_square ;
        END
    END B3
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.9300 0.6225 1.0350 0.7875 ;
        RECT 0.4650 0.7125 0.9300 0.7875 ;
        VIA 0.9825 0.6975 VIA12_square ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.2075 0.8625 1.3575 0.9375 ;
        RECT 1.2075 0.5625 1.3125 0.6375 ;
        RECT 1.1325 0.5625 1.2075 0.9375 ;
        RECT 0.6975 0.8625 1.1325 0.9375 ;
        VIA 1.2300 0.6000 VIA12_square ;
        END
    END B1
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.6225 0.2625 1.0875 0.3375 ;
        RECT 0.6225 0.5325 0.6525 0.6375 ;
        RECT 0.5475 0.2625 0.6225 0.6375 ;
        VIA 0.5850 0.5325 VIA12_square ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.3450 0.8625 0.5775 0.9375 ;
        RECT 0.2400 0.7350 0.3450 0.9375 ;
        RECT 0.0600 0.8625 0.2400 0.9375 ;
        VIA 0.2925 0.8175 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1500 0.4650 0.2400 0.5850 ;
        RECT 0.1425 0.4650 0.1500 0.6825 ;
        RECT 0.0375 0.3675 0.1425 0.6825 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.8450 -0.0750 1.8900 0.0750 ;
        RECT 1.7250 -0.0750 1.8450 0.2175 ;
        RECT 1.4250 -0.0750 1.7250 0.0750 ;
        RECT 1.3050 -0.0750 1.4250 0.1800 ;
        RECT 1.0050 -0.0750 1.3050 0.0750 ;
        RECT 0.8850 -0.0750 1.0050 0.1800 ;
        RECT 0.0000 -0.0750 0.8850 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.8450 0.9750 1.8900 1.1250 ;
        RECT 1.7250 0.8175 1.8450 1.1250 ;
        RECT 1.4250 0.9750 1.7250 1.1250 ;
        RECT 1.3050 0.8700 1.4250 1.1250 ;
        RECT 0.1650 0.9750 1.3050 1.1250 ;
        RECT 0.0450 0.7875 0.1650 1.1250 ;
        RECT 0.0000 0.9750 0.0450 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.7550 0.1575 1.8150 0.2175 ;
        RECT 1.7550 0.8325 1.8150 0.8925 ;
        RECT 1.6425 0.4950 1.7025 0.5550 ;
        RECT 1.5450 0.2775 1.6050 0.3375 ;
        RECT 1.5450 0.7650 1.6050 0.8250 ;
        RECT 1.4400 0.4950 1.5000 0.5550 ;
        RECT 1.3350 0.1200 1.3950 0.1800 ;
        RECT 1.3350 0.8700 1.3950 0.9300 ;
        RECT 1.2300 0.4950 1.2900 0.5550 ;
        RECT 1.1250 0.2400 1.1850 0.3000 ;
        RECT 1.0125 0.4950 1.0725 0.5550 ;
        RECT 0.9150 0.1200 0.9750 0.1800 ;
        RECT 0.8100 0.4950 0.8700 0.5550 ;
        RECT 0.7050 0.3150 0.7650 0.3750 ;
        RECT 0.7050 0.8325 0.7650 0.8925 ;
        RECT 0.5925 0.4950 0.6525 0.5550 ;
        RECT 0.4950 0.1650 0.5550 0.2250 ;
        RECT 0.3900 0.4950 0.4500 0.5550 ;
        RECT 0.2850 0.3150 0.3450 0.3750 ;
        RECT 0.1800 0.4950 0.2400 0.5550 ;
        RECT 0.0750 0.1875 0.1350 0.2475 ;
        RECT 0.0750 0.8175 0.1350 0.8775 ;
        LAYER M1 ;
        RECT 1.4625 0.4650 1.7025 0.5850 ;
        RECT 1.3875 0.2550 1.4625 0.7950 ;
        RECT 1.2975 0.2550 1.3875 0.3375 ;
        RECT 1.2300 0.7200 1.3875 0.7950 ;
        RECT 1.1475 0.4500 1.3125 0.6450 ;
        RECT 1.1550 0.7200 1.2300 0.9000 ;
        RECT 1.1025 0.2100 1.1925 0.3300 ;
        RECT 0.6750 0.8250 1.1550 0.9000 ;
        RECT 0.8400 0.2550 1.1025 0.3300 ;
        RECT 0.9975 0.4350 1.0725 0.7500 ;
        RECT 0.8775 0.6450 0.9975 0.7500 ;
        RECT 0.8025 0.4650 0.9225 0.5700 ;
        RECT 0.7650 0.2550 0.8400 0.3825 ;
        RECT 0.7275 0.4650 0.8025 0.7200 ;
        RECT 0.2550 0.3075 0.7650 0.3825 ;
        RECT 0.5325 0.4575 0.6525 0.7350 ;
        RECT 0.1500 0.1575 0.5850 0.2325 ;
        RECT 0.3225 0.4650 0.4575 0.9000 ;
        RECT 0.2400 0.7350 0.3225 0.9000 ;
        RECT 0.0450 0.1575 0.1500 0.2775 ;
        LAYER VIA1 ;
        RECT 1.3425 0.2550 1.4175 0.3300 ;
        RECT 0.3825 0.1575 0.4575 0.2325 ;
        LAYER M2 ;
        RECT 1.3200 0.2550 1.4625 0.3300 ;
        RECT 1.2450 0.1125 1.3200 0.3300 ;
        RECT 0.4725 0.1125 1.2450 0.1875 ;
        RECT 0.3675 0.1125 0.4725 0.2700 ;
    END
END OA33_0011


MACRO OA33_0111
    CLASS CORE ;
    FOREIGN OA33_0111 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.7800 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 3.0975 0.2400 3.4125 0.7500 ;
        VIA 3.2550 0.3225 VIA12_slot ;
        VIA 3.2550 0.6675 VIA12_slot ;
        END
    END Z
    PIN B3
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.6825 0.2625 0.7875 0.6075 ;
        RECT 0.2100 0.2625 0.6825 0.3375 ;
        VIA 0.7350 0.5250 VIA12_square ;
        END
    END B3
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.6075 0.7125 1.0575 0.7875 ;
        RECT 0.5025 0.6075 0.6075 0.7875 ;
        VIA 0.5550 0.6900 VIA12_square ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.1775 0.4725 1.2825 0.9375 ;
        RECT 0.4275 0.8625 1.1775 0.9375 ;
        RECT 0.3525 0.5625 0.4275 0.9375 ;
        RECT 0.1425 0.5625 0.3525 0.6375 ;
        VIA 1.2300 0.5550 VIA12_square ;
        VIA 0.2250 0.6000 VIA12_square ;
        END
    END B1
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.9425 0.2625 2.0475 0.6075 ;
        RECT 1.4700 0.2625 1.9425 0.3375 ;
        VIA 1.9950 0.5250 VIA12_square ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.8075 0.7125 2.2725 0.7875 ;
        RECT 1.7325 0.6075 1.8075 0.7875 ;
        VIA 1.7700 0.6900 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 2.4450 0.4350 2.5500 0.9375 ;
        RECT 1.5825 0.8625 2.4450 0.9375 ;
        RECT 1.4775 0.4725 1.5825 0.9375 ;
        VIA 2.4975 0.5250 VIA12_square ;
        VIA 1.5300 0.5550 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 3.7125 -0.0750 3.7800 0.0750 ;
        RECT 3.6375 -0.0750 3.7125 0.3150 ;
        RECT 3.3150 -0.0750 3.6375 0.0750 ;
        RECT 3.1950 -0.0750 3.3150 0.1950 ;
        RECT 2.8950 -0.0750 3.1950 0.0750 ;
        RECT 2.7900 -0.0750 2.8950 0.2475 ;
        RECT 1.2150 -0.0750 2.7900 0.0750 ;
        RECT 1.0950 -0.0750 1.2150 0.2025 ;
        RECT 0.7950 -0.0750 1.0950 0.0750 ;
        RECT 0.6750 -0.0750 0.7950 0.2025 ;
        RECT 0.3750 -0.0750 0.6750 0.0750 ;
        RECT 0.2550 -0.0750 0.3750 0.2025 ;
        RECT 0.0000 -0.0750 0.2550 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 3.7125 0.9750 3.7800 1.1250 ;
        RECT 3.6375 0.6375 3.7125 1.1250 ;
        RECT 3.3075 0.9750 3.6375 1.1250 ;
        RECT 3.2025 0.8025 3.3075 1.1250 ;
        RECT 2.8950 0.9750 3.2025 1.1250 ;
        RECT 2.7750 0.8025 2.8950 1.1250 ;
        RECT 2.6850 0.9750 2.7750 1.1250 ;
        RECT 2.5650 0.8025 2.6850 1.1250 ;
        RECT 1.4250 0.9750 2.5650 1.1250 ;
        RECT 1.3050 0.8625 1.4250 1.1250 ;
        RECT 0.1650 0.9750 1.3050 1.1250 ;
        RECT 0.0450 0.7650 0.1650 1.1250 ;
        RECT 0.0000 0.9750 0.0450 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 3.6450 0.2250 3.7050 0.2850 ;
        RECT 3.6450 0.6675 3.7050 0.7275 ;
        RECT 3.6450 0.8325 3.7050 0.8925 ;
        RECT 3.5400 0.4650 3.6000 0.5250 ;
        RECT 3.4350 0.2250 3.4950 0.2850 ;
        RECT 3.4350 0.7575 3.4950 0.8175 ;
        RECT 3.3300 0.4650 3.3900 0.5250 ;
        RECT 3.2250 0.1275 3.2850 0.1875 ;
        RECT 3.2250 0.8325 3.2850 0.8925 ;
        RECT 3.1200 0.4650 3.1800 0.5250 ;
        RECT 3.0150 0.2250 3.0750 0.2850 ;
        RECT 3.0150 0.7575 3.0750 0.8175 ;
        RECT 2.9100 0.4650 2.9700 0.5250 ;
        RECT 2.8050 0.1575 2.8650 0.2175 ;
        RECT 2.8050 0.8100 2.8650 0.8700 ;
        RECT 2.5950 0.1725 2.6550 0.2325 ;
        RECT 2.5950 0.8100 2.6550 0.8700 ;
        RECT 2.4900 0.4950 2.5500 0.5550 ;
        RECT 2.3850 0.3225 2.4450 0.3825 ;
        RECT 2.2800 0.4950 2.3400 0.5550 ;
        RECT 2.1750 0.1725 2.2350 0.2325 ;
        RECT 2.0700 0.4950 2.1300 0.5550 ;
        RECT 1.9650 0.3225 2.0250 0.3825 ;
        RECT 1.9650 0.8175 2.0250 0.8775 ;
        RECT 1.8600 0.4950 1.9200 0.5550 ;
        RECT 1.7550 0.1725 1.8150 0.2325 ;
        RECT 1.6500 0.4950 1.7100 0.5550 ;
        RECT 1.5450 0.3225 1.6050 0.3825 ;
        RECT 1.4400 0.4950 1.5000 0.5550 ;
        RECT 1.3350 0.2325 1.3950 0.2925 ;
        RECT 1.3350 0.8700 1.3950 0.9300 ;
        RECT 1.2300 0.4950 1.2900 0.5550 ;
        RECT 1.1250 0.1350 1.1850 0.1950 ;
        RECT 1.0200 0.4950 1.0800 0.5550 ;
        RECT 0.9150 0.2850 0.9750 0.3450 ;
        RECT 0.8100 0.4950 0.8700 0.5550 ;
        RECT 0.7050 0.1350 0.7650 0.1950 ;
        RECT 0.7050 0.8175 0.7650 0.8775 ;
        RECT 0.6000 0.4950 0.6600 0.5550 ;
        RECT 0.4950 0.2850 0.5550 0.3450 ;
        RECT 0.3900 0.4950 0.4500 0.5550 ;
        RECT 0.2850 0.1350 0.3450 0.1950 ;
        RECT 0.1800 0.4650 0.2400 0.5250 ;
        RECT 0.0750 0.2625 0.1350 0.3225 ;
        RECT 0.0750 0.8325 0.1350 0.8925 ;
        LAYER M1 ;
        RECT 2.9100 0.4425 3.6300 0.5475 ;
        RECT 3.4125 0.1950 3.5175 0.3675 ;
        RECT 3.4275 0.6225 3.5025 0.8700 ;
        RECT 3.0825 0.6225 3.4275 0.7125 ;
        RECT 3.0975 0.2775 3.4125 0.3675 ;
        RECT 2.9925 0.1950 3.0975 0.3675 ;
        RECT 3.0075 0.6225 3.0825 0.8700 ;
        RECT 2.8350 0.3225 2.9100 0.7275 ;
        RECT 2.6775 0.3225 2.8350 0.3975 ;
        RECT 2.4900 0.6525 2.8350 0.7275 ;
        RECT 2.4225 0.4725 2.7225 0.5775 ;
        RECT 1.4025 0.1650 2.6850 0.2400 ;
        RECT 2.6100 0.3150 2.6775 0.3975 ;
        RECT 1.5075 0.3150 2.6100 0.3900 ;
        RECT 2.4150 0.6525 2.4900 0.8850 ;
        RECT 1.5750 0.8100 2.4150 0.8850 ;
        RECT 2.2350 0.4650 2.3400 0.7275 ;
        RECT 1.7550 0.6525 2.2350 0.7275 ;
        RECT 1.8300 0.4725 2.1600 0.5775 ;
        RECT 1.6500 0.4650 1.7550 0.7275 ;
        RECT 1.3800 0.4725 1.5750 0.6375 ;
        RECT 1.5000 0.7125 1.5750 0.8850 ;
        RECT 1.2300 0.7125 1.5000 0.7875 ;
        RECT 1.3275 0.1650 1.4025 0.3525 ;
        RECT 0.1425 0.2775 1.3275 0.3525 ;
        RECT 1.1550 0.4275 1.3050 0.6375 ;
        RECT 1.1550 0.7125 1.2300 0.8850 ;
        RECT 0.6675 0.8100 1.1550 0.8850 ;
        RECT 0.9750 0.4650 1.0800 0.7275 ;
        RECT 0.4950 0.6525 0.9750 0.7275 ;
        RECT 0.5700 0.4725 0.9000 0.5775 ;
        RECT 0.3825 0.4650 0.4950 0.7275 ;
        RECT 0.1125 0.4275 0.3075 0.6375 ;
        RECT 0.0675 0.2325 0.1425 0.3525 ;
    END
END OA33_0111


MACRO OA33_1000
    CLASS CORE ;
    FOREIGN OA33_1000 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.6800 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 1.5675 0.1500 1.6425 0.9000 ;
        RECT 1.5375 0.1500 1.5675 0.3825 ;
        RECT 1.5375 0.6675 1.5675 0.9000 ;
        END
    END Z
    PIN B3
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.8625 0.4125 1.3200 0.4875 ;
        RECT 0.7575 0.4125 0.8625 0.5850 ;
        VIA 0.8100 0.5025 VIA12_square ;
        END
    END B3
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.9300 0.6225 1.0350 0.7875 ;
        RECT 0.4650 0.7125 0.9300 0.7875 ;
        VIA 0.9825 0.6975 VIA12_square ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.2075 0.8625 1.3575 0.9375 ;
        RECT 1.2075 0.5625 1.3125 0.6375 ;
        RECT 1.1325 0.5625 1.2075 0.9375 ;
        RECT 0.6975 0.8625 1.1325 0.9375 ;
        VIA 1.2300 0.6000 VIA12_square ;
        END
    END B1
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.6225 0.2625 1.0875 0.3375 ;
        RECT 0.6225 0.5325 0.6525 0.6375 ;
        RECT 0.5475 0.2625 0.6225 0.6375 ;
        VIA 0.5850 0.5325 VIA12_square ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.3450 0.8625 0.5775 0.9375 ;
        RECT 0.2400 0.7350 0.3450 0.9375 ;
        RECT 0.0600 0.8625 0.2400 0.9375 ;
        VIA 0.2925 0.8175 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1500 0.4650 0.2400 0.5850 ;
        RECT 0.1425 0.4650 0.1500 0.6825 ;
        RECT 0.0375 0.3675 0.1425 0.6825 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.4250 -0.0750 1.6800 0.0750 ;
        RECT 1.3050 -0.0750 1.4250 0.1800 ;
        RECT 1.0050 -0.0750 1.3050 0.0750 ;
        RECT 0.8850 -0.0750 1.0050 0.1800 ;
        RECT 0.0000 -0.0750 0.8850 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.4250 0.9750 1.6800 1.1250 ;
        RECT 1.3050 0.8700 1.4250 1.1250 ;
        RECT 0.1650 0.9750 1.3050 1.1250 ;
        RECT 0.0450 0.7875 0.1650 1.1250 ;
        RECT 0.0000 0.9750 0.0450 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.5450 0.1800 1.6050 0.2400 ;
        RECT 1.5450 0.8100 1.6050 0.8700 ;
        RECT 1.4325 0.4950 1.4925 0.5550 ;
        RECT 1.3350 0.1200 1.3950 0.1800 ;
        RECT 1.3350 0.8700 1.3950 0.9300 ;
        RECT 1.2300 0.4950 1.2900 0.5550 ;
        RECT 1.1250 0.1800 1.1850 0.2400 ;
        RECT 1.0125 0.4950 1.0725 0.5550 ;
        RECT 0.9150 0.1200 0.9750 0.1800 ;
        RECT 0.8100 0.4950 0.8700 0.5550 ;
        RECT 0.7050 0.3150 0.7650 0.3750 ;
        RECT 0.7050 0.8325 0.7650 0.8925 ;
        RECT 0.5925 0.4950 0.6525 0.5550 ;
        RECT 0.4950 0.1650 0.5550 0.2250 ;
        RECT 0.3900 0.4950 0.4500 0.5550 ;
        RECT 0.2850 0.3150 0.3450 0.3750 ;
        RECT 0.1800 0.4950 0.2400 0.5550 ;
        RECT 0.0750 0.1875 0.1350 0.2475 ;
        RECT 0.0750 0.8175 0.1350 0.8775 ;
        LAYER M1 ;
        RECT 1.4625 0.4650 1.4925 0.5850 ;
        RECT 1.3875 0.2550 1.4625 0.7950 ;
        RECT 1.2975 0.2550 1.3875 0.3375 ;
        RECT 1.2300 0.7200 1.3875 0.7950 ;
        RECT 1.1475 0.4500 1.3125 0.6450 ;
        RECT 1.1550 0.7200 1.2300 0.9000 ;
        RECT 1.0875 0.1500 1.1925 0.3300 ;
        RECT 0.6750 0.8250 1.1550 0.9000 ;
        RECT 0.8400 0.2550 1.0875 0.3300 ;
        RECT 0.9975 0.4350 1.0725 0.7500 ;
        RECT 0.8775 0.6450 0.9975 0.7500 ;
        RECT 0.8025 0.4650 0.9225 0.5700 ;
        RECT 0.7650 0.2550 0.8400 0.3825 ;
        RECT 0.7275 0.4650 0.8025 0.7200 ;
        RECT 0.2550 0.3075 0.7650 0.3825 ;
        RECT 0.5325 0.4575 0.6525 0.7350 ;
        RECT 0.1500 0.1575 0.5850 0.2325 ;
        RECT 0.3225 0.4650 0.4575 0.9000 ;
        RECT 0.2400 0.7350 0.3225 0.9000 ;
        RECT 0.0450 0.1575 0.1500 0.2775 ;
        LAYER VIA1 ;
        RECT 1.3425 0.2550 1.4175 0.3300 ;
        RECT 0.3825 0.1575 0.4575 0.2325 ;
        LAYER M2 ;
        RECT 1.3200 0.2550 1.4625 0.3300 ;
        RECT 1.2450 0.1125 1.3200 0.3300 ;
        RECT 0.4725 0.1125 1.2450 0.1875 ;
        RECT 0.3675 0.1125 0.4725 0.2700 ;
    END
END OA33_1000


MACRO OA33_1010
    CLASS CORE ;
    FOREIGN OA33_1010 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.6800 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 1.5675 0.2175 1.6425 0.8325 ;
        RECT 1.5375 0.2175 1.5675 0.3825 ;
        RECT 1.5375 0.6675 1.5675 0.8325 ;
        END
    END Z
    PIN B3
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.8625 0.4125 1.3200 0.4875 ;
        RECT 0.7575 0.4125 0.8625 0.5850 ;
        VIA 0.8100 0.5025 VIA12_square ;
        END
    END B3
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.9300 0.6225 1.0350 0.7875 ;
        RECT 0.4650 0.7125 0.9300 0.7875 ;
        VIA 0.9825 0.6975 VIA12_square ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.2075 0.8625 1.3575 0.9375 ;
        RECT 1.2075 0.5625 1.3125 0.6375 ;
        RECT 1.1325 0.5625 1.2075 0.9375 ;
        RECT 0.6975 0.8625 1.1325 0.9375 ;
        VIA 1.2300 0.6000 VIA12_square ;
        END
    END B1
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.6225 0.2625 1.0875 0.3375 ;
        RECT 0.6225 0.5325 0.6525 0.6375 ;
        RECT 0.5475 0.2625 0.6225 0.6375 ;
        VIA 0.5850 0.5325 VIA12_square ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.3450 0.8625 0.5775 0.9375 ;
        RECT 0.2400 0.7350 0.3450 0.9375 ;
        RECT 0.0600 0.8625 0.2400 0.9375 ;
        VIA 0.2925 0.8175 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1500 0.4650 0.2400 0.5850 ;
        RECT 0.1425 0.4650 0.1500 0.6825 ;
        RECT 0.0375 0.3675 0.1425 0.6825 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.4250 -0.0750 1.6800 0.0750 ;
        RECT 1.3050 -0.0750 1.4250 0.1800 ;
        RECT 1.0050 -0.0750 1.3050 0.0750 ;
        RECT 0.8850 -0.0750 1.0050 0.1800 ;
        RECT 0.0000 -0.0750 0.8850 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.4250 0.9750 1.6800 1.1250 ;
        RECT 1.3050 0.8700 1.4250 1.1250 ;
        RECT 0.1650 0.9750 1.3050 1.1250 ;
        RECT 0.0450 0.7875 0.1650 1.1250 ;
        RECT 0.0000 0.9750 0.0450 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.5450 0.2700 1.6050 0.3300 ;
        RECT 1.5450 0.7200 1.6050 0.7800 ;
        RECT 1.4325 0.4950 1.4925 0.5550 ;
        RECT 1.3350 0.1200 1.3950 0.1800 ;
        RECT 1.3350 0.8700 1.3950 0.9300 ;
        RECT 1.2300 0.4950 1.2900 0.5550 ;
        RECT 1.1250 0.2400 1.1850 0.3000 ;
        RECT 1.0125 0.4950 1.0725 0.5550 ;
        RECT 0.9150 0.1200 0.9750 0.1800 ;
        RECT 0.8100 0.4950 0.8700 0.5550 ;
        RECT 0.7050 0.3150 0.7650 0.3750 ;
        RECT 0.7050 0.8325 0.7650 0.8925 ;
        RECT 0.5925 0.4950 0.6525 0.5550 ;
        RECT 0.4950 0.1650 0.5550 0.2250 ;
        RECT 0.3900 0.4950 0.4500 0.5550 ;
        RECT 0.2850 0.3150 0.3450 0.3750 ;
        RECT 0.1800 0.4950 0.2400 0.5550 ;
        RECT 0.0750 0.1875 0.1350 0.2475 ;
        RECT 0.0750 0.8175 0.1350 0.8775 ;
        LAYER M1 ;
        RECT 1.4625 0.4650 1.4925 0.5850 ;
        RECT 1.3875 0.2550 1.4625 0.7950 ;
        RECT 1.2975 0.2550 1.3875 0.3375 ;
        RECT 1.2300 0.7200 1.3875 0.7950 ;
        RECT 1.1475 0.4500 1.3125 0.6450 ;
        RECT 1.1550 0.7200 1.2300 0.9000 ;
        RECT 1.1025 0.2100 1.1925 0.3300 ;
        RECT 0.6750 0.8250 1.1550 0.9000 ;
        RECT 0.8400 0.2550 1.1025 0.3300 ;
        RECT 0.9975 0.4350 1.0725 0.7500 ;
        RECT 0.8775 0.6450 0.9975 0.7500 ;
        RECT 0.8025 0.4650 0.9225 0.5700 ;
        RECT 0.7650 0.2550 0.8400 0.3825 ;
        RECT 0.7275 0.4650 0.8025 0.7200 ;
        RECT 0.2550 0.3075 0.7650 0.3825 ;
        RECT 0.5325 0.4575 0.6525 0.7350 ;
        RECT 0.1500 0.1575 0.5850 0.2325 ;
        RECT 0.3225 0.4650 0.4575 0.9000 ;
        RECT 0.2400 0.7350 0.3225 0.9000 ;
        RECT 0.0450 0.1575 0.1500 0.2775 ;
        LAYER VIA1 ;
        RECT 1.3425 0.2550 1.4175 0.3300 ;
        RECT 0.3825 0.1575 0.4575 0.2325 ;
        LAYER M2 ;
        RECT 1.3200 0.2550 1.4625 0.3300 ;
        RECT 1.2450 0.1125 1.3200 0.3300 ;
        RECT 0.4725 0.1125 1.2450 0.1875 ;
        RECT 0.3675 0.1125 0.4725 0.2700 ;
    END
END OA33_1010


MACRO OAI211_0011
    CLASS CORE ;
    FOREIGN OAI211_0011 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.8900 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 0.8175 0.7125 1.3875 0.7875 ;
        RECT 0.7725 0.2625 0.8175 0.7875 ;
        RECT 0.7125 0.2625 0.7725 0.9300 ;
        RECT 0.6675 0.7125 0.7125 0.9300 ;
        VIA 1.2750 0.7500 VIA12_square ;
        VIA 0.7650 0.3375 VIA12_square ;
        VIA 0.7200 0.8475 VIA12_square ;
        END
    END ZN
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.9600 0.4125 1.4250 0.4875 ;
        VIA 1.3125 0.4500 VIA12_square ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.9600 0.5625 1.7700 0.6375 ;
        VIA 1.6575 0.6000 VIA12_square ;
        VIA 1.0725 0.6000 VIA12_square ;
        END
    END B
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.5625 0.1125 1.0275 0.1875 ;
        RECT 0.5625 0.4500 0.5925 0.6000 ;
        RECT 0.4875 0.1125 0.5625 0.6000 ;
        VIA 0.5400 0.5250 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.8175 0.4575 0.8925 0.5700 ;
        RECT 0.7425 0.4575 0.8175 0.7350 ;
        RECT 0.2925 0.6600 0.7425 0.7350 ;
        RECT 0.2175 0.4875 0.2925 0.7350 ;
        RECT 0.1425 0.4875 0.2175 0.6825 ;
        RECT 0.0675 0.3675 0.1425 0.6825 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.4250 -0.0750 1.8900 0.0750 ;
        RECT 1.3050 -0.0750 1.4250 0.1875 ;
        RECT 0.0000 -0.0750 1.3050 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.8225 0.9750 1.8900 1.1250 ;
        RECT 1.7475 0.7425 1.8225 1.1250 ;
        RECT 1.4250 0.9750 1.7475 1.1250 ;
        RECT 1.3050 0.8625 1.4250 1.1250 ;
        RECT 0.9825 0.9750 1.3050 1.1250 ;
        RECT 0.9075 0.7875 0.9825 1.1250 ;
        RECT 0.1425 0.9750 0.9075 1.1250 ;
        RECT 0.0675 0.7875 0.1425 1.1250 ;
        RECT 0.0000 0.9750 0.0675 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.7550 0.2250 1.8150 0.2850 ;
        RECT 1.7550 0.7725 1.8150 0.8325 ;
        RECT 1.6500 0.4950 1.7100 0.5550 ;
        RECT 1.5450 0.7575 1.6050 0.8175 ;
        RECT 1.4400 0.4950 1.5000 0.5550 ;
        RECT 1.3350 0.1275 1.3950 0.1875 ;
        RECT 1.3350 0.8625 1.3950 0.9225 ;
        RECT 1.2300 0.4950 1.2900 0.5550 ;
        RECT 1.1250 0.7575 1.1850 0.8175 ;
        RECT 1.0200 0.4725 1.0800 0.5325 ;
        RECT 0.9150 0.1575 0.9750 0.2175 ;
        RECT 0.9150 0.8175 0.9750 0.8775 ;
        RECT 0.8100 0.4875 0.8700 0.5475 ;
        RECT 0.7050 0.3075 0.7650 0.3675 ;
        RECT 0.6000 0.4950 0.6600 0.5550 ;
        RECT 0.4950 0.1575 0.5550 0.2175 ;
        RECT 0.4950 0.8175 0.5550 0.8775 ;
        RECT 0.3900 0.4950 0.4500 0.5550 ;
        RECT 0.2850 0.3075 0.3450 0.3675 ;
        RECT 0.1800 0.4950 0.2400 0.5550 ;
        RECT 0.0750 0.1800 0.1350 0.2400 ;
        RECT 0.0750 0.8175 0.1350 0.8775 ;
        LAYER M1 ;
        RECT 1.7400 0.1875 1.8300 0.3375 ;
        RECT 1.5750 0.4725 1.7850 0.6375 ;
        RECT 1.2150 0.2625 1.7400 0.3375 ;
        RECT 1.5300 0.7125 1.6200 0.8550 ;
        RECT 1.2150 0.7125 1.5300 0.7875 ;
        RECT 1.2300 0.4125 1.5000 0.5850 ;
        RECT 1.1400 0.1500 1.2150 0.3375 ;
        RECT 1.0950 0.7125 1.2150 0.8400 ;
        RECT 0.9675 0.4200 1.1550 0.6375 ;
        RECT 0.1575 0.1500 1.1400 0.2250 ;
        RECT 0.2550 0.3000 0.8625 0.3825 ;
        RECT 0.3675 0.8100 0.8025 0.9000 ;
        RECT 0.3825 0.4650 0.6675 0.5850 ;
        RECT 0.0525 0.1500 0.1575 0.2625 ;
    END
END OAI211_0011


MACRO OAI211_0100
    CLASS CORE ;
    FOREIGN OAI211_0100 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.2400 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 4.0350 0.2850 4.1925 0.4050 ;
        RECT 4.0350 0.6375 4.1925 0.7575 ;
        RECT 3.7200 0.2850 4.0350 0.7575 ;
        RECT 3.5625 0.2850 3.7200 0.4050 ;
        RECT 3.5625 0.6375 3.7200 0.7575 ;
        VIA 4.0350 0.3450 VIA12_slot ;
        VIA 4.0350 0.6975 VIA12_slot ;
        VIA 3.7200 0.3450 VIA12_slot ;
        VIA 3.7200 0.6975 VIA12_slot ;
        END
    END ZN
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 9.0975 0.4050 9.1725 0.6900 ;
        RECT 9.0075 0.4050 9.0975 0.5700 ;
        RECT 6.6600 0.4650 9.0075 0.5700 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 4.7250 0.4125 5.0850 0.4875 ;
        RECT 4.6200 0.4125 4.7250 0.6375 ;
        VIA 4.6725 0.5250 VIA12_square ;
        END
    END B
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 2.7450 0.4500 2.8500 0.6375 ;
        RECT 2.3250 0.5625 2.7450 0.6375 ;
        VIA 2.7975 0.5325 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.3225 0.4650 2.5725 0.5700 ;
        RECT 0.1425 0.4650 0.3225 0.6450 ;
        RECT 0.0675 0.3675 0.1425 0.6450 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 8.9850 -0.0750 9.2400 0.0750 ;
        RECT 8.8650 -0.0750 8.9850 0.1800 ;
        RECT 8.5650 -0.0750 8.8650 0.0750 ;
        RECT 8.4450 -0.0750 8.5650 0.1800 ;
        RECT 8.1450 -0.0750 8.4450 0.0750 ;
        RECT 8.0250 -0.0750 8.1450 0.1800 ;
        RECT 7.7250 -0.0750 8.0250 0.0750 ;
        RECT 7.6050 -0.0750 7.7250 0.1800 ;
        RECT 7.3050 -0.0750 7.6050 0.0750 ;
        RECT 7.1850 -0.0750 7.3050 0.1800 ;
        RECT 6.8850 -0.0750 7.1850 0.0750 ;
        RECT 6.7650 -0.0750 6.8850 0.1800 ;
        RECT 0.0000 -0.0750 6.7650 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 9.1875 0.9750 9.2400 1.1250 ;
        RECT 9.0825 0.8100 9.1875 1.1250 ;
        RECT 8.7750 0.9750 9.0825 1.1250 ;
        RECT 8.6550 0.8325 8.7750 1.1250 ;
        RECT 8.3550 0.9750 8.6550 1.1250 ;
        RECT 8.2350 0.8325 8.3550 1.1250 ;
        RECT 7.9350 0.9750 8.2350 1.1250 ;
        RECT 7.8150 0.8325 7.9350 1.1250 ;
        RECT 7.5150 0.9750 7.8150 1.1250 ;
        RECT 7.3950 0.8325 7.5150 1.1250 ;
        RECT 7.0950 0.9750 7.3950 1.1250 ;
        RECT 6.9750 0.8325 7.0950 1.1250 ;
        RECT 6.6750 0.9750 6.9750 1.1250 ;
        RECT 6.5550 0.8325 6.6750 1.1250 ;
        RECT 6.2550 0.9750 6.5550 1.1250 ;
        RECT 6.1350 0.8325 6.2550 1.1250 ;
        RECT 5.8350 0.9750 6.1350 1.1250 ;
        RECT 5.7150 0.8325 5.8350 1.1250 ;
        RECT 5.4150 0.9750 5.7150 1.1250 ;
        RECT 5.2950 0.8325 5.4150 1.1250 ;
        RECT 4.9950 0.9750 5.2950 1.1250 ;
        RECT 4.8750 0.8700 4.9950 1.1250 ;
        RECT 4.5750 0.9750 4.8750 1.1250 ;
        RECT 4.4550 0.8325 4.5750 1.1250 ;
        RECT 2.4750 0.9750 4.4550 1.1250 ;
        RECT 2.3550 0.8700 2.4750 1.1250 ;
        RECT 2.0550 0.9750 2.3550 1.1250 ;
        RECT 1.9350 0.8700 2.0550 1.1250 ;
        RECT 1.6350 0.9750 1.9350 1.1250 ;
        RECT 1.5150 0.8700 1.6350 1.1250 ;
        RECT 1.2150 0.9750 1.5150 1.1250 ;
        RECT 1.0950 0.8700 1.2150 1.1250 ;
        RECT 0.7950 0.9750 1.0950 1.1250 ;
        RECT 0.6750 0.8700 0.7950 1.1250 ;
        RECT 0.3750 0.9750 0.6750 1.1250 ;
        RECT 0.2550 0.8700 0.3750 1.1250 ;
        RECT 0.0000 0.9750 0.2550 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 9.1050 0.2400 9.1650 0.3000 ;
        RECT 9.1050 0.8325 9.1650 0.8925 ;
        RECT 9.0000 0.4950 9.0600 0.5550 ;
        RECT 8.8950 0.1200 8.9550 0.1800 ;
        RECT 8.8950 0.7500 8.9550 0.8100 ;
        RECT 8.7900 0.4950 8.8500 0.5550 ;
        RECT 8.6850 0.2850 8.7450 0.3450 ;
        RECT 8.6850 0.8325 8.7450 0.8925 ;
        RECT 8.5800 0.4950 8.6400 0.5550 ;
        RECT 8.4750 0.1200 8.5350 0.1800 ;
        RECT 8.4750 0.7500 8.5350 0.8100 ;
        RECT 8.3700 0.4950 8.4300 0.5550 ;
        RECT 8.2650 0.3075 8.3250 0.3675 ;
        RECT 8.2650 0.8325 8.3250 0.8925 ;
        RECT 8.1600 0.4950 8.2200 0.5550 ;
        RECT 8.0550 0.1200 8.1150 0.1800 ;
        RECT 8.0550 0.7500 8.1150 0.8100 ;
        RECT 7.9500 0.4950 8.0100 0.5550 ;
        RECT 7.8450 0.3075 7.9050 0.3675 ;
        RECT 7.8450 0.8325 7.9050 0.8925 ;
        RECT 7.7400 0.4950 7.8000 0.5550 ;
        RECT 7.6350 0.1200 7.6950 0.1800 ;
        RECT 7.6350 0.7500 7.6950 0.8100 ;
        RECT 7.5300 0.4950 7.5900 0.5550 ;
        RECT 7.4250 0.3075 7.4850 0.3675 ;
        RECT 7.4250 0.8325 7.4850 0.8925 ;
        RECT 7.3200 0.4950 7.3800 0.5550 ;
        RECT 7.2150 0.1200 7.2750 0.1800 ;
        RECT 7.2150 0.7500 7.2750 0.8100 ;
        RECT 7.1100 0.4950 7.1700 0.5550 ;
        RECT 7.0050 0.3075 7.0650 0.3675 ;
        RECT 7.0050 0.8325 7.0650 0.8925 ;
        RECT 6.9000 0.4950 6.9600 0.5550 ;
        RECT 6.7950 0.1200 6.8550 0.1800 ;
        RECT 6.7950 0.7500 6.8550 0.8100 ;
        RECT 6.6900 0.4950 6.7500 0.5550 ;
        RECT 6.5850 0.3075 6.6450 0.3675 ;
        RECT 6.5850 0.8325 6.6450 0.8925 ;
        RECT 6.3750 0.1575 6.4350 0.2175 ;
        RECT 6.2700 0.4950 6.3300 0.5550 ;
        RECT 6.1650 0.3075 6.2250 0.3675 ;
        RECT 6.1650 0.8325 6.2250 0.8925 ;
        RECT 6.0600 0.4950 6.1200 0.5550 ;
        RECT 5.9550 0.1575 6.0150 0.2175 ;
        RECT 5.9550 0.7500 6.0150 0.8100 ;
        RECT 5.8500 0.4950 5.9100 0.5550 ;
        RECT 5.7450 0.3075 5.8050 0.3675 ;
        RECT 5.7450 0.8325 5.8050 0.8925 ;
        RECT 5.6400 0.4950 5.7000 0.5550 ;
        RECT 5.5350 0.1575 5.5950 0.2175 ;
        RECT 5.5350 0.7500 5.5950 0.8100 ;
        RECT 5.4300 0.4950 5.4900 0.5550 ;
        RECT 5.3250 0.3075 5.3850 0.3675 ;
        RECT 5.3250 0.8325 5.3850 0.8925 ;
        RECT 5.2200 0.4950 5.2800 0.5550 ;
        RECT 5.1150 0.1575 5.1750 0.2175 ;
        RECT 5.1150 0.7500 5.1750 0.8100 ;
        RECT 5.0100 0.4950 5.0700 0.5550 ;
        RECT 4.9050 0.3075 4.9650 0.3675 ;
        RECT 4.9050 0.8700 4.9650 0.9300 ;
        RECT 4.8000 0.4950 4.8600 0.5550 ;
        RECT 4.6950 0.1575 4.7550 0.2175 ;
        RECT 4.6950 0.7275 4.7550 0.7875 ;
        RECT 4.5900 0.4950 4.6500 0.5550 ;
        RECT 4.4850 0.3075 4.5450 0.3675 ;
        RECT 4.4850 0.8325 4.5450 0.8925 ;
        RECT 4.3800 0.4950 4.4400 0.5550 ;
        RECT 4.2750 0.1575 4.3350 0.2175 ;
        RECT 4.2750 0.8175 4.3350 0.8775 ;
        RECT 4.1625 0.4950 4.2225 0.5550 ;
        RECT 4.0650 0.3075 4.1250 0.3675 ;
        RECT 4.0650 0.6900 4.1250 0.7500 ;
        RECT 3.9600 0.4950 4.0200 0.5550 ;
        RECT 3.8550 0.1575 3.9150 0.2175 ;
        RECT 3.8550 0.8325 3.9150 0.8925 ;
        RECT 3.7500 0.4950 3.8100 0.5550 ;
        RECT 3.6450 0.3075 3.7050 0.3675 ;
        RECT 3.6450 0.6900 3.7050 0.7500 ;
        RECT 3.5400 0.4950 3.6000 0.5550 ;
        RECT 3.4350 0.1575 3.4950 0.2175 ;
        RECT 3.4350 0.8325 3.4950 0.8925 ;
        RECT 3.3300 0.4950 3.3900 0.5550 ;
        RECT 3.2250 0.3075 3.2850 0.3675 ;
        RECT 3.2250 0.6900 3.2850 0.7500 ;
        RECT 3.1200 0.4950 3.1800 0.5550 ;
        RECT 3.0150 0.1575 3.0750 0.2175 ;
        RECT 3.0150 0.8325 3.0750 0.8925 ;
        RECT 2.9100 0.4950 2.9700 0.5550 ;
        RECT 2.8050 0.3075 2.8650 0.3675 ;
        RECT 2.8050 0.6900 2.8650 0.7500 ;
        RECT 2.7000 0.4950 2.7600 0.5550 ;
        RECT 2.5950 0.1575 2.6550 0.2175 ;
        RECT 2.5950 0.7575 2.6550 0.8175 ;
        RECT 2.4900 0.4875 2.5500 0.5475 ;
        RECT 2.3850 0.3075 2.4450 0.3675 ;
        RECT 2.3850 0.8700 2.4450 0.9300 ;
        RECT 2.2800 0.4875 2.3400 0.5475 ;
        RECT 2.1750 0.1575 2.2350 0.2175 ;
        RECT 2.1750 0.7275 2.2350 0.7875 ;
        RECT 2.0700 0.4875 2.1300 0.5475 ;
        RECT 1.9650 0.3075 2.0250 0.3675 ;
        RECT 1.9650 0.8700 2.0250 0.9300 ;
        RECT 1.8600 0.4875 1.9200 0.5475 ;
        RECT 1.7550 0.1575 1.8150 0.2175 ;
        RECT 1.7550 0.7275 1.8150 0.7875 ;
        RECT 1.6500 0.4875 1.7100 0.5475 ;
        RECT 1.5450 0.8700 1.6050 0.9300 ;
        RECT 1.4400 0.4875 1.5000 0.5475 ;
        RECT 1.3350 0.1575 1.3950 0.2175 ;
        RECT 1.3350 0.7275 1.3950 0.7875 ;
        RECT 1.2300 0.4875 1.2900 0.5475 ;
        RECT 1.1250 0.3075 1.1850 0.3675 ;
        RECT 1.1250 0.8700 1.1850 0.9300 ;
        RECT 1.0200 0.4875 1.0800 0.5475 ;
        RECT 0.9150 0.1575 0.9750 0.2175 ;
        RECT 0.9150 0.7275 0.9750 0.7875 ;
        RECT 0.8100 0.4875 0.8700 0.5475 ;
        RECT 0.7050 0.8700 0.7650 0.9300 ;
        RECT 0.6000 0.4875 0.6600 0.5475 ;
        RECT 0.4950 0.1575 0.5550 0.2175 ;
        RECT 0.4950 0.7275 0.5550 0.7875 ;
        RECT 0.3900 0.4875 0.4500 0.5475 ;
        RECT 0.2850 0.3075 0.3450 0.3675 ;
        RECT 0.2850 0.8700 0.3450 0.9300 ;
        RECT 0.1800 0.4875 0.2400 0.5475 ;
        RECT 0.0750 0.1725 0.1350 0.2325 ;
        RECT 0.0750 0.7575 0.1350 0.8175 ;
        LAYER M1 ;
        RECT 9.0975 0.2100 9.1725 0.3300 ;
        RECT 8.7525 0.2550 9.0975 0.3300 ;
        RECT 8.8875 0.6450 8.9625 0.8475 ;
        RECT 8.5425 0.6450 8.8875 0.7575 ;
        RECT 8.6775 0.2550 8.7525 0.3750 ;
        RECT 4.4400 0.3000 8.6775 0.3750 ;
        RECT 8.4675 0.6450 8.5425 0.8475 ;
        RECT 8.1225 0.6450 8.4675 0.7575 ;
        RECT 8.0475 0.6450 8.1225 0.8475 ;
        RECT 7.7025 0.6450 8.0475 0.7575 ;
        RECT 7.6275 0.6450 7.7025 0.8475 ;
        RECT 7.2825 0.6450 7.6275 0.7575 ;
        RECT 7.2075 0.6450 7.2825 0.8475 ;
        RECT 6.8625 0.6450 7.2075 0.7575 ;
        RECT 6.7875 0.6450 6.8625 0.8475 ;
        RECT 6.0225 0.6450 6.7875 0.7575 ;
        RECT 0.1575 0.1500 6.4800 0.2250 ;
        RECT 4.3500 0.4650 6.3600 0.5700 ;
        RECT 5.9475 0.6450 6.0225 0.8475 ;
        RECT 5.6025 0.6450 5.9475 0.7575 ;
        RECT 5.5275 0.6450 5.6025 0.8475 ;
        RECT 5.1825 0.6450 5.5275 0.7575 ;
        RECT 5.1075 0.6450 5.1825 0.8475 ;
        RECT 4.7625 0.6450 5.1075 0.7575 ;
        RECT 4.6875 0.6450 4.7625 0.8475 ;
        RECT 4.4175 0.6450 4.6875 0.7500 ;
        RECT 4.1775 0.6450 4.4175 0.7200 ;
        RECT 4.2525 0.7950 4.3575 0.9000 ;
        RECT 2.6550 0.4650 4.2525 0.5700 ;
        RECT 2.6625 0.8250 4.2525 0.9000 ;
        RECT 0.2475 0.3000 4.1925 0.3900 ;
        RECT 2.7750 0.6450 4.1775 0.7500 ;
        RECT 2.5875 0.7200 2.6625 0.9000 ;
        RECT 0.1425 0.7200 2.5875 0.7950 ;
        RECT 0.0525 0.1500 0.1575 0.2550 ;
        RECT 0.0675 0.7200 0.1425 0.8475 ;
        LAYER M2 ;
        RECT 4.0650 0.2850 4.1925 0.4050 ;
        RECT 4.0650 0.6375 4.1925 0.7575 ;
        RECT 3.5625 0.2850 3.6900 0.4050 ;
        RECT 3.5625 0.6375 3.6900 0.7575 ;
    END
END OAI211_0100


MACRO OAI211_0111
    CLASS CORE ;
    FOREIGN OAI211_0111 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.7800 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 1.2075 0.2700 1.5225 0.7800 ;
        VIA 1.3650 0.3525 VIA12_slot ;
        VIA 1.3650 0.6975 VIA12_slot ;
        END
    END ZN
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 3.2925 0.4125 3.5700 0.4875 ;
        RECT 3.2175 0.4125 3.2925 0.6375 ;
        RECT 2.9400 0.5625 3.2175 0.6375 ;
        VIA 3.2550 0.5325 VIA12_square ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 2.6625 0.4125 2.9400 0.4875 ;
        RECT 2.5875 0.4125 2.6625 0.6375 ;
        RECT 2.3100 0.5625 2.5875 0.6375 ;
        VIA 2.6250 0.5325 VIA12_square ;
        END
    END B
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.6575 0.4125 2.1225 0.4875 ;
        VIA 1.7850 0.4500 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.5625 0.4125 0.8400 0.4875 ;
        RECT 0.4875 0.4125 0.5625 0.6375 ;
        RECT 0.2100 0.5625 0.4875 0.6375 ;
        VIA 0.5250 0.5325 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 3.5175 -0.0750 3.7800 0.0750 ;
        RECT 3.4125 -0.0750 3.5175 0.2250 ;
        RECT 3.0975 -0.0750 3.4125 0.0750 ;
        RECT 2.9925 -0.0750 3.0975 0.2250 ;
        RECT 0.0000 -0.0750 2.9925 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 3.5175 0.9750 3.7800 1.1250 ;
        RECT 3.4125 0.8325 3.5175 1.1250 ;
        RECT 3.0975 0.9750 3.4125 1.1250 ;
        RECT 2.9925 0.8325 3.0975 1.1250 ;
        RECT 2.6775 0.9750 2.9925 1.1250 ;
        RECT 2.5725 0.8325 2.6775 1.1250 ;
        RECT 2.2575 0.9750 2.5725 1.1250 ;
        RECT 2.1525 0.8325 2.2575 1.1250 ;
        RECT 0.7950 0.9750 2.1525 1.1250 ;
        RECT 0.6750 0.8325 0.7950 1.1250 ;
        RECT 0.3750 0.9750 0.6750 1.1250 ;
        RECT 0.2550 0.8325 0.3750 1.1250 ;
        RECT 0.0000 0.9750 0.2550 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 3.6450 0.2925 3.7050 0.3525 ;
        RECT 3.6450 0.6825 3.7050 0.7425 ;
        RECT 3.5400 0.4950 3.6000 0.5550 ;
        RECT 3.4350 0.1425 3.4950 0.2025 ;
        RECT 3.4350 0.8550 3.4950 0.9150 ;
        RECT 3.3300 0.4950 3.3900 0.5550 ;
        RECT 3.2250 0.3075 3.2850 0.3675 ;
        RECT 3.2250 0.6675 3.2850 0.7275 ;
        RECT 3.1200 0.4950 3.1800 0.5550 ;
        RECT 3.0150 0.1425 3.0750 0.2025 ;
        RECT 3.0150 0.8550 3.0750 0.9150 ;
        RECT 2.9100 0.4950 2.9700 0.5550 ;
        RECT 2.8050 0.3075 2.8650 0.3675 ;
        RECT 2.8050 0.6675 2.8650 0.7275 ;
        RECT 2.7000 0.4950 2.7600 0.5550 ;
        RECT 2.5950 0.1575 2.6550 0.2175 ;
        RECT 2.5950 0.8550 2.6550 0.9150 ;
        RECT 2.4900 0.4950 2.5500 0.5550 ;
        RECT 2.3850 0.3075 2.4450 0.3675 ;
        RECT 2.3850 0.6675 2.4450 0.7275 ;
        RECT 2.2800 0.4950 2.3400 0.5550 ;
        RECT 2.1750 0.1575 2.2350 0.2175 ;
        RECT 2.1750 0.8550 2.2350 0.9150 ;
        RECT 2.0700 0.4950 2.1300 0.5550 ;
        RECT 1.9650 0.3075 2.0250 0.3675 ;
        RECT 1.9650 0.6825 2.0250 0.7425 ;
        RECT 1.7550 0.1575 1.8150 0.2175 ;
        RECT 1.7550 0.8325 1.8150 0.8925 ;
        RECT 1.6500 0.4950 1.7100 0.5550 ;
        RECT 1.5450 0.3225 1.6050 0.3825 ;
        RECT 1.5450 0.6675 1.6050 0.7275 ;
        RECT 1.4400 0.4950 1.5000 0.5550 ;
        RECT 1.3350 0.1575 1.3950 0.2175 ;
        RECT 1.3350 0.8325 1.3950 0.8925 ;
        RECT 1.2300 0.4950 1.2900 0.5550 ;
        RECT 1.1250 0.3150 1.1850 0.3750 ;
        RECT 1.1250 0.6825 1.1850 0.7425 ;
        RECT 1.0275 0.4950 1.0875 0.5550 ;
        RECT 0.9150 0.1575 0.9750 0.2175 ;
        RECT 0.9150 0.8325 0.9750 0.8925 ;
        RECT 0.8100 0.4950 0.8700 0.5550 ;
        RECT 0.7050 0.3225 0.7650 0.3825 ;
        RECT 0.7050 0.8400 0.7650 0.9000 ;
        RECT 0.6000 0.4950 0.6600 0.5550 ;
        RECT 0.4950 0.1575 0.5550 0.2175 ;
        RECT 0.4950 0.6900 0.5550 0.7500 ;
        RECT 0.3900 0.4950 0.4500 0.5550 ;
        RECT 0.2850 0.3225 0.3450 0.3825 ;
        RECT 0.2850 0.8400 0.3450 0.9000 ;
        RECT 0.0750 0.1950 0.1350 0.2550 ;
        RECT 0.0750 0.7275 0.1350 0.7875 ;
        RECT 0.1800 0.4950 0.2400 0.5550 ;
        LAYER M1 ;
        RECT 1.2225 0.6450 3.7350 0.7500 ;
        RECT 3.6225 0.2700 3.7275 0.3750 ;
        RECT 2.8725 0.4650 3.6300 0.5700 ;
        RECT 1.9350 0.3000 3.6225 0.3750 ;
        RECT 2.0325 0.4650 2.7900 0.5700 ;
        RECT 0.1575 0.1500 2.6850 0.2250 ;
        RECT 0.9450 0.8250 1.8450 0.9000 ;
        RECT 1.7475 0.3300 1.8225 0.5700 ;
        RECT 1.1025 0.4800 1.7475 0.5700 ;
        RECT 0.2625 0.3000 1.6275 0.4050 ;
        RECT 1.0950 0.6750 1.2225 0.7500 ;
        RECT 0.9975 0.4800 1.1025 0.5850 ;
        RECT 0.8700 0.6825 0.9450 0.9000 ;
        RECT 0.1350 0.4800 0.9000 0.5850 ;
        RECT 0.1575 0.6825 0.8700 0.7575 ;
        RECT 0.0525 0.1500 0.1575 0.2775 ;
        RECT 0.0525 0.6825 0.1575 0.8175 ;
    END
END OAI211_0111


MACRO OAI211_1000
    CLASS CORE ;
    FOREIGN OAI211_1000 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.0500 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 0.6075 0.6825 0.6975 0.7875 ;
        RECT 0.5325 0.2625 0.6075 0.7875 ;
        RECT 0.4725 0.2625 0.5325 0.4275 ;
        RECT 0.0675 0.2625 0.4725 0.3375 ;
        VIA 0.6150 0.7425 VIA12_square ;
        VIA 0.5100 0.3450 VIA12_square ;
        END
    END ZN
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.9075 0.3675 0.9825 0.6825 ;
        RECT 0.8175 0.4800 0.9075 0.6000 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.8175 0.1125 0.9825 0.1875 ;
        RECT 0.7125 0.1125 0.8175 0.3150 ;
        RECT 0.4125 0.1125 0.7125 0.1875 ;
        VIA 0.7650 0.2325 VIA12_square ;
        END
    END B
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1425 0.4800 0.2325 0.6000 ;
        RECT 0.0675 0.3675 0.1425 0.6825 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.4275 0.8625 0.6075 0.9375 ;
        RECT 0.3525 0.5100 0.4275 0.9375 ;
        RECT 0.0675 0.8625 0.3525 0.9375 ;
        VIA 0.3900 0.5925 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.0125 -0.0750 1.0500 0.0750 ;
        RECT 0.9075 -0.0750 1.0125 0.2475 ;
        RECT 0.0000 -0.0750 0.9075 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.9975 0.9750 1.0500 1.1250 ;
        RECT 0.8925 0.8100 0.9975 1.1250 ;
        RECT 0.5850 0.9750 0.8925 1.1250 ;
        RECT 0.4650 0.8700 0.5850 1.1250 ;
        RECT 0.0000 0.9750 0.4650 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 0.9150 0.1575 0.9750 0.2175 ;
        RECT 0.9150 0.8325 0.9750 0.8925 ;
        RECT 0.8175 0.5100 0.8775 0.5700 ;
        RECT 0.7050 0.7800 0.7650 0.8400 ;
        RECT 0.6000 0.5100 0.6600 0.5700 ;
        RECT 0.4950 0.1575 0.5550 0.2175 ;
        RECT 0.4950 0.8700 0.5550 0.9300 ;
        RECT 0.3900 0.5100 0.4500 0.5700 ;
        RECT 0.2850 0.3075 0.3450 0.3675 ;
        RECT 0.1725 0.5100 0.2325 0.5700 ;
        RECT 0.0750 0.1800 0.1350 0.2400 ;
        RECT 0.0750 0.8175 0.1350 0.8775 ;
        LAYER M1 ;
        RECT 0.7425 0.1500 0.8175 0.4050 ;
        RECT 0.6825 0.7050 0.7950 0.8700 ;
        RECT 0.7125 0.1500 0.7425 0.6000 ;
        RECT 0.6675 0.3300 0.7125 0.6000 ;
        RECT 0.3825 0.7050 0.6825 0.7800 ;
        RECT 0.6000 0.4800 0.6675 0.6000 ;
        RECT 0.2550 0.3000 0.5925 0.4050 ;
        RECT 0.1425 0.1500 0.5850 0.2250 ;
        RECT 0.3075 0.4800 0.5250 0.6300 ;
        RECT 0.3075 0.7050 0.3825 0.9000 ;
        RECT 0.0525 0.7950 0.3075 0.9000 ;
        RECT 0.0675 0.1500 0.1425 0.2700 ;
    END
END OAI211_1000


MACRO OAI211_1010
    CLASS CORE ;
    FOREIGN OAI211_1010 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.2600 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 1.1025 0.7200 1.2075 0.8400 ;
        RECT 0.6675 0.7200 1.1025 0.7950 ;
        RECT 0.5925 0.3000 0.6675 0.7950 ;
        RECT 0.2550 0.3000 0.5925 0.3750 ;
        RECT 0.4800 0.6750 0.5925 0.7950 ;
        END
    END ZN
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.0200 0.4125 1.1850 0.6375 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.7575 0.4125 0.9225 0.6375 ;
        END
    END B
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.3900 0.4500 0.4500 0.5700 ;
        RECT 0.3150 0.4500 0.3900 0.8325 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1425 0.4500 0.2400 0.5700 ;
        RECT 0.0675 0.3675 0.1425 0.6825 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.2150 -0.0750 1.2600 0.0750 ;
        RECT 1.0950 -0.0750 1.2150 0.2925 ;
        RECT 0.0000 -0.0750 1.0950 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.0050 0.9750 1.2600 1.1250 ;
        RECT 0.8850 0.8700 1.0050 1.1250 ;
        RECT 0.1650 0.9750 0.8850 1.1250 ;
        RECT 0.0450 0.8025 0.1650 1.1250 ;
        RECT 0.0000 0.9750 0.0450 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.1250 0.2250 1.1850 0.2850 ;
        RECT 1.1250 0.7500 1.1850 0.8100 ;
        RECT 1.0200 0.4800 1.0800 0.5400 ;
        RECT 0.9150 0.8700 0.9750 0.9300 ;
        RECT 0.8100 0.4800 0.8700 0.5400 ;
        RECT 0.7050 0.1575 0.7650 0.2175 ;
        RECT 0.7050 0.7275 0.7650 0.7875 ;
        RECT 0.4950 0.1575 0.5550 0.2175 ;
        RECT 0.4950 0.7050 0.5550 0.7650 ;
        RECT 0.3900 0.4800 0.4500 0.5400 ;
        RECT 0.2850 0.3075 0.3450 0.3675 ;
        RECT 0.1800 0.4800 0.2400 0.5400 ;
        RECT 0.0750 0.1725 0.1350 0.2325 ;
        RECT 0.0750 0.8100 0.1350 0.8700 ;
        LAYER M1 ;
        RECT 0.1575 0.1500 0.7950 0.2250 ;
        RECT 0.0525 0.1500 0.1575 0.2550 ;
    END
END OAI211_1010


MACRO OAI21_0011
    CLASS CORE ;
    FOREIGN OAI21_0011 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.4700 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 0.8925 0.8625 1.2075 0.9375 ;
        RECT 0.8175 0.2625 0.8925 0.9375 ;
        RECT 0.7875 0.2625 0.8175 0.4200 ;
        RECT 0.3525 0.7125 0.8175 0.7875 ;
        VIA 0.8550 0.8550 VIA12_square ;
        VIA 0.8400 0.3375 VIA12_square ;
        VIA 0.5100 0.7500 VIA12_square ;
        END
    END ZN
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1425 0.4125 0.4800 0.5325 ;
        RECT 0.0675 0.4125 0.1425 0.6825 ;
        END
    END B
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.6075 0.2625 0.7125 0.5775 ;
        RECT 0.2100 0.2625 0.6075 0.3375 ;
        VIA 0.6600 0.5025 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.9825 0.1125 1.0875 0.6000 ;
        RECT 0.5475 0.1125 0.9825 0.1875 ;
        VIA 1.0350 0.5175 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.3750 -0.0750 1.4700 0.0750 ;
        RECT 0.2550 -0.0750 0.3750 0.1800 ;
        RECT 0.0000 -0.0750 0.2550 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.4175 0.9750 1.4700 1.1250 ;
        RECT 1.3125 0.8025 1.4175 1.1250 ;
        RECT 0.5850 0.9750 1.3125 1.1250 ;
        RECT 0.4650 0.8625 0.5850 1.1250 ;
        RECT 0.1425 0.9750 0.4650 1.1250 ;
        RECT 0.0675 0.7875 0.1425 1.1250 ;
        RECT 0.0000 0.9750 0.0675 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.3350 0.1800 1.3950 0.2400 ;
        RECT 1.3350 0.8325 1.3950 0.8925 ;
        RECT 1.2300 0.4950 1.2900 0.5550 ;
        RECT 1.1250 0.3075 1.1850 0.3675 ;
        RECT 1.0200 0.4875 1.0800 0.5475 ;
        RECT 0.9150 0.1575 0.9750 0.2175 ;
        RECT 0.9150 0.8175 0.9750 0.8775 ;
        RECT 0.8175 0.4875 0.8775 0.5475 ;
        RECT 0.7050 0.3075 0.7650 0.3675 ;
        RECT 0.6000 0.4875 0.6600 0.5475 ;
        RECT 0.4950 0.2100 0.5550 0.2700 ;
        RECT 0.4950 0.8625 0.5550 0.9225 ;
        RECT 0.3900 0.4650 0.4500 0.5250 ;
        RECT 0.2850 0.1200 0.3450 0.1800 ;
        RECT 0.2850 0.7050 0.3450 0.7650 ;
        RECT 0.1800 0.4650 0.2400 0.5250 ;
        RECT 0.0750 0.2400 0.1350 0.3000 ;
        RECT 0.0750 0.8325 0.1350 0.8925 ;
        LAYER M1 ;
        RECT 1.3350 0.1500 1.4100 0.2850 ;
        RECT 0.5550 0.1500 1.3350 0.2250 ;
        RECT 1.2750 0.4875 1.3275 0.5625 ;
        RECT 1.2000 0.4875 1.2750 0.7350 ;
        RECT 0.6750 0.3000 1.2300 0.3750 ;
        RECT 0.7200 0.8100 1.2075 0.9000 ;
        RECT 0.7425 0.6600 1.2000 0.7350 ;
        RECT 0.8175 0.4500 1.1250 0.5850 ;
        RECT 0.6675 0.4500 0.7425 0.7350 ;
        RECT 0.5775 0.4500 0.6675 0.5775 ;
        RECT 0.2550 0.6825 0.5925 0.7875 ;
        RECT 0.4800 0.1500 0.5550 0.3300 ;
        RECT 0.1575 0.2550 0.4800 0.3300 ;
        RECT 0.0675 0.2100 0.1575 0.3300 ;
    END
END OAI21_0011


MACRO OAI21_0100
    CLASS CORE ;
    FOREIGN OAI21_0100 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.1400 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 3.6225 0.2850 3.7800 0.4050 ;
        RECT 3.6225 0.6300 3.7800 0.7500 ;
        RECT 3.3075 0.2850 3.6225 0.7500 ;
        RECT 3.1500 0.2850 3.3075 0.4050 ;
        RECT 3.1500 0.6300 3.3075 0.7500 ;
        VIA 3.6225 0.3450 VIA12_slot ;
        VIA 3.6225 0.6900 VIA12_slot ;
        VIA 3.3075 0.3450 VIA12_slot ;
        VIA 3.3075 0.6900 VIA12_slot ;
        END
    END ZN
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 6.9375 0.4125 7.1025 0.6375 ;
        RECT 4.5600 0.4650 6.9375 0.5700 ;
        END
    END B
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.2025 0.5625 0.6675 0.6375 ;
        VIA 0.3150 0.6000 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 4.4400 0.5625 4.8225 0.6375 ;
        RECT 4.3350 0.4275 4.4400 0.6375 ;
        VIA 4.3875 0.5175 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 6.8850 -0.0750 7.1400 0.0750 ;
        RECT 6.7650 -0.0750 6.8850 0.1875 ;
        RECT 6.4650 -0.0750 6.7650 0.0750 ;
        RECT 6.3450 -0.0750 6.4650 0.2325 ;
        RECT 6.0450 -0.0750 6.3450 0.0750 ;
        RECT 5.9250 -0.0750 6.0450 0.2325 ;
        RECT 5.6250 -0.0750 5.9250 0.0750 ;
        RECT 5.5050 -0.0750 5.6250 0.2325 ;
        RECT 5.2050 -0.0750 5.5050 0.0750 ;
        RECT 5.0850 -0.0750 5.2050 0.2325 ;
        RECT 4.7850 -0.0750 5.0850 0.0750 ;
        RECT 4.6650 -0.0750 4.7850 0.2325 ;
        RECT 0.0000 -0.0750 4.6650 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 7.0725 0.9750 7.1400 1.1250 ;
        RECT 6.9975 0.7875 7.0725 1.1250 ;
        RECT 6.6675 0.9750 6.9975 1.1250 ;
        RECT 6.5625 0.8100 6.6675 1.1250 ;
        RECT 6.2475 0.9750 6.5625 1.1250 ;
        RECT 6.1425 0.8100 6.2475 1.1250 ;
        RECT 5.8275 0.9750 6.1425 1.1250 ;
        RECT 5.7225 0.8100 5.8275 1.1250 ;
        RECT 5.4075 0.9750 5.7225 1.1250 ;
        RECT 5.3025 0.8100 5.4075 1.1250 ;
        RECT 4.9875 0.9750 5.3025 1.1250 ;
        RECT 4.8825 0.8100 4.9875 1.1250 ;
        RECT 4.5750 0.9750 4.8825 1.1250 ;
        RECT 4.4700 0.8025 4.5750 1.1250 ;
        RECT 2.4675 0.9750 4.4700 1.1250 ;
        RECT 2.3625 0.8250 2.4675 1.1250 ;
        RECT 2.0475 0.9750 2.3625 1.1250 ;
        RECT 1.9425 0.8250 2.0475 1.1250 ;
        RECT 1.6275 0.9750 1.9425 1.1250 ;
        RECT 1.5225 0.8250 1.6275 1.1250 ;
        RECT 1.2075 0.9750 1.5225 1.1250 ;
        RECT 1.1025 0.8250 1.2075 1.1250 ;
        RECT 0.7875 0.9750 1.1025 1.1250 ;
        RECT 0.6825 0.8250 0.7875 1.1250 ;
        RECT 0.3750 0.9750 0.6825 1.1250 ;
        RECT 0.2550 0.8625 0.3750 1.1250 ;
        RECT 0.0000 0.9750 0.2550 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 7.0050 0.2250 7.0650 0.2850 ;
        RECT 7.0050 0.8325 7.0650 0.8925 ;
        RECT 6.9000 0.4950 6.9600 0.5550 ;
        RECT 6.7950 0.1275 6.8550 0.1875 ;
        RECT 6.7950 0.8100 6.8550 0.8700 ;
        RECT 6.6900 0.4950 6.7500 0.5550 ;
        RECT 6.5850 0.3150 6.6450 0.3750 ;
        RECT 6.5850 0.8325 6.6450 0.8925 ;
        RECT 6.4800 0.4950 6.5400 0.5550 ;
        RECT 6.3750 0.1425 6.4350 0.2025 ;
        RECT 6.3750 0.8100 6.4350 0.8700 ;
        RECT 6.2700 0.4950 6.3300 0.5550 ;
        RECT 6.1650 0.3150 6.2250 0.3750 ;
        RECT 6.1650 0.8325 6.2250 0.8925 ;
        RECT 6.0600 0.4950 6.1200 0.5550 ;
        RECT 5.9550 0.1425 6.0150 0.2025 ;
        RECT 5.9550 0.8100 6.0150 0.8700 ;
        RECT 5.8500 0.4950 5.9100 0.5550 ;
        RECT 5.7450 0.3150 5.8050 0.3750 ;
        RECT 5.7450 0.8325 5.8050 0.8925 ;
        RECT 5.6400 0.4875 5.7000 0.5475 ;
        RECT 5.5350 0.1425 5.5950 0.2025 ;
        RECT 5.5350 0.8100 5.5950 0.8700 ;
        RECT 5.4300 0.4875 5.4900 0.5475 ;
        RECT 5.3250 0.3150 5.3850 0.3750 ;
        RECT 5.3250 0.8325 5.3850 0.8925 ;
        RECT 5.2200 0.4875 5.2800 0.5475 ;
        RECT 5.1150 0.1425 5.1750 0.2025 ;
        RECT 5.1150 0.8100 5.1750 0.8700 ;
        RECT 5.0100 0.4875 5.0700 0.5475 ;
        RECT 4.9050 0.3150 4.9650 0.3750 ;
        RECT 4.9050 0.8325 4.9650 0.8925 ;
        RECT 4.8000 0.4875 4.8600 0.5475 ;
        RECT 4.6950 0.1425 4.7550 0.2025 ;
        RECT 4.6950 0.6675 4.7550 0.7275 ;
        RECT 4.5900 0.4875 4.6500 0.5475 ;
        RECT 4.4850 0.2175 4.5450 0.2775 ;
        RECT 4.4850 0.8325 4.5450 0.8925 ;
        RECT 4.2750 0.3075 4.3350 0.3675 ;
        RECT 4.2750 0.8325 4.3350 0.8925 ;
        RECT 4.1700 0.4950 4.2300 0.5550 ;
        RECT 4.0650 0.1575 4.1250 0.2175 ;
        RECT 4.0650 0.6675 4.1250 0.7275 ;
        RECT 3.9600 0.4950 4.0200 0.5550 ;
        RECT 3.8550 0.3150 3.9150 0.3750 ;
        RECT 3.8550 0.8325 3.9150 0.8925 ;
        RECT 3.7500 0.4950 3.8100 0.5550 ;
        RECT 3.6450 0.1575 3.7050 0.2175 ;
        RECT 3.6450 0.6675 3.7050 0.7275 ;
        RECT 3.5400 0.4950 3.6000 0.5550 ;
        RECT 3.4350 0.3150 3.4950 0.3750 ;
        RECT 3.4350 0.8325 3.4950 0.8925 ;
        RECT 3.3300 0.4950 3.3900 0.5550 ;
        RECT 3.2250 0.1575 3.2850 0.2175 ;
        RECT 3.2250 0.6675 3.2850 0.7275 ;
        RECT 3.1200 0.4950 3.1800 0.5550 ;
        RECT 3.0150 0.3150 3.0750 0.3750 ;
        RECT 3.0150 0.8325 3.0750 0.8925 ;
        RECT 2.9100 0.4950 2.9700 0.5550 ;
        RECT 2.8050 0.1575 2.8650 0.2175 ;
        RECT 2.8050 0.6675 2.8650 0.7275 ;
        RECT 2.7000 0.4950 2.7600 0.5550 ;
        RECT 2.5950 0.3150 2.6550 0.3750 ;
        RECT 2.5950 0.7575 2.6550 0.8175 ;
        RECT 2.4900 0.4950 2.5500 0.5550 ;
        RECT 2.3850 0.1575 2.4450 0.2175 ;
        RECT 2.3850 0.8475 2.4450 0.9075 ;
        RECT 2.2800 0.4950 2.3400 0.5550 ;
        RECT 2.1750 0.3150 2.2350 0.3750 ;
        RECT 2.1750 0.6825 2.2350 0.7425 ;
        RECT 2.0700 0.4950 2.1300 0.5550 ;
        RECT 1.9650 0.1575 2.0250 0.2175 ;
        RECT 1.9650 0.8475 2.0250 0.9075 ;
        RECT 1.8600 0.4950 1.9200 0.5550 ;
        RECT 1.7550 0.3150 1.8150 0.3750 ;
        RECT 1.7550 0.6825 1.8150 0.7425 ;
        RECT 1.6500 0.4950 1.7100 0.5550 ;
        RECT 1.5450 0.1575 1.6050 0.2175 ;
        RECT 1.5450 0.8475 1.6050 0.9075 ;
        RECT 1.4400 0.4950 1.5000 0.5550 ;
        RECT 1.3350 0.6825 1.3950 0.7425 ;
        RECT 1.2300 0.4950 1.2900 0.5550 ;
        RECT 1.1250 0.1575 1.1850 0.2175 ;
        RECT 1.1250 0.8475 1.1850 0.9075 ;
        RECT 1.0200 0.4950 1.0800 0.5550 ;
        RECT 0.9150 0.3150 0.9750 0.3750 ;
        RECT 0.9150 0.6825 0.9750 0.7425 ;
        RECT 0.8100 0.4950 0.8700 0.5550 ;
        RECT 0.7050 0.1575 0.7650 0.2175 ;
        RECT 0.7050 0.8475 0.7650 0.9075 ;
        RECT 0.6000 0.4950 0.6600 0.5550 ;
        RECT 0.4950 0.6975 0.5550 0.7575 ;
        RECT 0.3900 0.4950 0.4500 0.5550 ;
        RECT 0.2850 0.1575 0.3450 0.2175 ;
        RECT 0.2850 0.8625 0.3450 0.9225 ;
        RECT 0.1800 0.4950 0.2400 0.5550 ;
        RECT 0.0750 0.2550 0.1350 0.3150 ;
        RECT 0.0750 0.7575 0.1350 0.8175 ;
        LAYER M1 ;
        RECT 6.9975 0.1800 7.0725 0.3375 ;
        RECT 6.8625 0.2625 6.9975 0.3375 ;
        RECT 6.8475 0.7800 6.8775 0.9000 ;
        RECT 6.7875 0.2625 6.8625 0.3825 ;
        RECT 6.7725 0.6450 6.8475 0.9000 ;
        RECT 4.5525 0.3075 6.7875 0.3825 ;
        RECT 6.4575 0.6450 6.7725 0.7275 ;
        RECT 6.3525 0.6450 6.4575 0.9000 ;
        RECT 6.0375 0.6450 6.3525 0.7275 ;
        RECT 5.9325 0.6450 6.0375 0.9000 ;
        RECT 5.6175 0.6450 5.9325 0.7275 ;
        RECT 5.5125 0.6450 5.6175 0.9000 ;
        RECT 5.1975 0.6450 5.5125 0.7275 ;
        RECT 5.0925 0.6450 5.1975 0.9000 ;
        RECT 2.7750 0.6450 5.0925 0.7275 ;
        RECT 4.4775 0.1500 4.5525 0.3825 ;
        RECT 0.2475 0.1500 4.4775 0.2250 ;
        RECT 2.6700 0.4650 4.4700 0.5700 ;
        RECT 0.1425 0.3000 4.3725 0.3900 ;
        RECT 2.6625 0.8250 4.3650 0.9000 ;
        RECT 2.5875 0.6750 2.6625 0.9000 ;
        RECT 0.5775 0.6750 2.5875 0.7500 ;
        RECT 0.3975 0.4725 2.5725 0.5775 ;
        RECT 0.4725 0.6750 0.5775 0.7875 ;
        RECT 0.1425 0.7125 0.4725 0.7875 ;
        RECT 0.2325 0.4725 0.3975 0.6375 ;
        RECT 0.1350 0.4725 0.2325 0.5775 ;
        RECT 0.0675 0.2250 0.1425 0.3900 ;
        RECT 0.0675 0.7125 0.1425 0.8625 ;
        LAYER M2 ;
        RECT 3.6525 0.2850 3.7800 0.4050 ;
        RECT 3.6525 0.6300 3.7800 0.7500 ;
        RECT 3.1500 0.2850 3.2775 0.4050 ;
        RECT 3.1500 0.6300 3.2775 0.7500 ;
    END
END OAI21_0100


MACRO OAI21_0111
    CLASS CORE ;
    FOREIGN OAI21_0111 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.9400 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 0.9975 0.2625 1.3125 0.7800 ;
        VIA 1.1550 0.3450 VIA12_slot ;
        VIA 1.1550 0.6975 VIA12_slot ;
        END
    END ZN
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 2.2425 0.4125 2.5125 0.4875 ;
        RECT 2.1675 0.4125 2.2425 0.6375 ;
        RECT 1.9275 0.5625 2.1675 0.6375 ;
        VIA 2.2050 0.5175 VIA12_square ;
        END
    END B
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.5625 0.4125 0.8325 0.4875 ;
        RECT 0.4875 0.4125 0.5625 0.6375 ;
        RECT 0.2475 0.5625 0.4875 0.6375 ;
        VIA 0.5250 0.5250 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.5225 0.4125 1.8825 0.4875 ;
        RECT 1.4175 0.4125 1.5225 0.5925 ;
        VIA 1.4700 0.5175 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 2.6850 -0.0750 2.9400 0.0750 ;
        RECT 2.5650 -0.0750 2.6850 0.2250 ;
        RECT 2.2650 -0.0750 2.5650 0.0750 ;
        RECT 2.1450 -0.0750 2.2650 0.2250 ;
        RECT 0.0000 -0.0750 2.1450 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 2.8875 0.9750 2.9400 1.1250 ;
        RECT 2.7825 0.6450 2.8875 1.1250 ;
        RECT 2.4675 0.9750 2.7825 1.1250 ;
        RECT 2.3625 0.8025 2.4675 1.1250 ;
        RECT 2.0550 0.9750 2.3625 1.1250 ;
        RECT 1.9500 0.8025 2.0550 1.1250 ;
        RECT 0.7800 0.9750 1.9500 1.1250 ;
        RECT 0.6750 0.8175 0.7800 1.1250 ;
        RECT 0.3675 0.9750 0.6750 1.1250 ;
        RECT 0.2625 0.8175 0.3675 1.1250 ;
        RECT 0.0000 0.9750 0.2625 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 2.8050 0.2775 2.8650 0.3375 ;
        RECT 2.8050 0.6675 2.8650 0.7275 ;
        RECT 2.8050 0.8325 2.8650 0.8925 ;
        RECT 2.7000 0.4875 2.7600 0.5475 ;
        RECT 2.5950 0.1500 2.6550 0.2100 ;
        RECT 2.5950 0.7575 2.6550 0.8175 ;
        RECT 2.4900 0.4875 2.5500 0.5475 ;
        RECT 2.3850 0.3075 2.4450 0.3675 ;
        RECT 2.3850 0.8325 2.4450 0.8925 ;
        RECT 2.2800 0.4875 2.3400 0.5475 ;
        RECT 2.1750 0.1500 2.2350 0.2100 ;
        RECT 2.1750 0.6600 2.2350 0.7200 ;
        RECT 2.0700 0.4875 2.1300 0.5475 ;
        RECT 1.9650 0.2175 2.0250 0.2775 ;
        RECT 1.9650 0.8325 2.0250 0.8925 ;
        RECT 1.7550 0.3075 1.8150 0.3675 ;
        RECT 1.7550 0.8325 1.8150 0.8925 ;
        RECT 1.6500 0.4875 1.7100 0.5475 ;
        RECT 1.5450 0.1575 1.6050 0.2175 ;
        RECT 1.5450 0.6675 1.6050 0.7275 ;
        RECT 1.4400 0.4875 1.5000 0.5475 ;
        RECT 1.3350 0.3075 1.3950 0.3675 ;
        RECT 1.3350 0.8325 1.3950 0.8925 ;
        RECT 1.2300 0.4875 1.2900 0.5475 ;
        RECT 1.1250 0.1575 1.1850 0.2175 ;
        RECT 1.1250 0.6825 1.1850 0.7425 ;
        RECT 1.0200 0.4875 1.0800 0.5475 ;
        RECT 0.9150 0.3075 0.9750 0.3675 ;
        RECT 0.9150 0.8325 0.9750 0.8925 ;
        RECT 0.8100 0.4950 0.8700 0.5550 ;
        RECT 0.7050 0.1575 0.7650 0.2175 ;
        RECT 0.7050 0.8475 0.7650 0.9075 ;
        RECT 0.6000 0.4950 0.6600 0.5550 ;
        RECT 0.4950 0.3075 0.5550 0.3675 ;
        RECT 0.4950 0.6750 0.5550 0.7350 ;
        RECT 0.3900 0.4950 0.4500 0.5550 ;
        RECT 0.2850 0.1575 0.3450 0.2175 ;
        RECT 0.2850 0.8475 0.3450 0.9075 ;
        RECT 0.1800 0.4950 0.2400 0.5550 ;
        RECT 0.0750 0.2550 0.1350 0.3150 ;
        RECT 0.0750 0.7275 0.1350 0.7875 ;
        LAYER M1 ;
        RECT 2.7825 0.2400 2.8800 0.3750 ;
        RECT 2.0400 0.4650 2.7900 0.5700 ;
        RECT 2.0325 0.3000 2.7825 0.3750 ;
        RECT 2.5875 0.6450 2.6625 0.8550 ;
        RECT 1.2975 0.6450 2.5875 0.7275 ;
        RECT 1.9575 0.1500 2.0325 0.3750 ;
        RECT 0.2475 0.1500 1.9575 0.2250 ;
        RECT 0.1425 0.3000 1.8450 0.3900 ;
        RECT 0.9300 0.8250 1.8450 0.9000 ;
        RECT 0.9900 0.4650 1.7400 0.5700 ;
        RECT 1.0125 0.6450 1.2975 0.7500 ;
        RECT 0.8550 0.6675 0.9300 0.9000 ;
        RECT 0.1500 0.4725 0.9000 0.5775 ;
        RECT 0.1425 0.6675 0.8550 0.7425 ;
        RECT 0.0675 0.2250 0.1425 0.3900 ;
        RECT 0.0675 0.6675 0.1425 0.8325 ;
    END
END OAI21_0111


MACRO OAI21_1000
    CLASS CORE ;
    FOREIGN OAI21_1000 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.0500 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.7350 0.6675 0.7875 0.9000 ;
        RECT 0.6600 0.3000 0.7350 0.9000 ;
        RECT 0.2550 0.3000 0.6600 0.3750 ;
        RECT 0.4650 0.8250 0.6600 0.9000 ;
        END
    END ZN
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.9075 0.3675 0.9825 0.6825 ;
        RECT 0.8100 0.4500 0.9075 0.5700 ;
        END
    END B
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1500 0.4575 0.2625 0.5625 ;
        RECT 0.0450 0.3675 0.1500 0.6825 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.3675 0.4500 0.4725 0.7500 ;
        RECT 0.3525 0.6675 0.3675 0.7500 ;
        RECT 0.2775 0.6675 0.3525 0.8325 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.9825 -0.0750 1.0500 0.0750 ;
        RECT 0.9075 -0.0750 0.9825 0.2475 ;
        RECT 0.0000 -0.0750 0.9075 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.9900 0.9750 1.0500 1.1250 ;
        RECT 0.9000 0.7875 0.9900 1.1250 ;
        RECT 0.1650 0.9750 0.9000 1.1250 ;
        RECT 0.0450 0.8175 0.1650 1.1250 ;
        RECT 0.0000 0.9750 0.0450 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 0.9150 0.1575 0.9750 0.2175 ;
        RECT 0.9150 0.8175 0.9750 0.8775 ;
        RECT 0.8100 0.4800 0.8700 0.5400 ;
        RECT 0.7050 0.1575 0.7650 0.2175 ;
        RECT 0.7050 0.8175 0.7650 0.8775 ;
        RECT 0.4950 0.1575 0.5550 0.2175 ;
        RECT 0.4950 0.8325 0.5550 0.8925 ;
        RECT 0.3900 0.4800 0.4500 0.5400 ;
        RECT 0.2850 0.3075 0.3450 0.3675 ;
        RECT 0.1800 0.4800 0.2400 0.5400 ;
        RECT 0.0750 0.1725 0.1350 0.2325 ;
        RECT 0.0750 0.8325 0.1350 0.8925 ;
        LAYER M1 ;
        RECT 0.1575 0.1500 0.7950 0.2250 ;
        RECT 0.0525 0.1500 0.1575 0.2550 ;
    END
END OAI21_1000


MACRO OAI21_1010
    CLASS CORE ;
    FOREIGN OAI21_1010 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.0500 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.7350 0.6675 0.7725 0.9000 ;
        RECT 0.6600 0.3000 0.7350 0.9000 ;
        RECT 0.2550 0.3000 0.6600 0.3750 ;
        RECT 0.4650 0.8250 0.6600 0.9000 ;
        END
    END ZN
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.9075 0.3675 0.9825 0.6825 ;
        RECT 0.8100 0.4500 0.9075 0.5700 ;
        END
    END B
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1500 0.4575 0.2625 0.5625 ;
        RECT 0.0450 0.3675 0.1500 0.6825 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.3675 0.4500 0.4725 0.7500 ;
        RECT 0.3525 0.6675 0.3675 0.7500 ;
        RECT 0.2775 0.6675 0.3525 0.8325 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.9825 -0.0750 1.0500 0.0750 ;
        RECT 0.9075 -0.0750 0.9825 0.2625 ;
        RECT 0.0000 -0.0750 0.9075 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.9900 0.9750 1.0500 1.1250 ;
        RECT 0.9000 0.7875 0.9900 1.1250 ;
        RECT 0.1650 0.9750 0.9000 1.1250 ;
        RECT 0.0450 0.7725 0.1650 1.1250 ;
        RECT 0.0000 0.9750 0.0450 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 0.9150 0.1725 0.9750 0.2325 ;
        RECT 0.9150 0.8175 0.9750 0.8775 ;
        RECT 0.8100 0.4800 0.8700 0.5400 ;
        RECT 0.7050 0.1575 0.7650 0.2175 ;
        RECT 0.7050 0.7500 0.7650 0.8100 ;
        RECT 0.4950 0.1575 0.5550 0.2175 ;
        RECT 0.4950 0.8325 0.5550 0.8925 ;
        RECT 0.3900 0.4800 0.4500 0.5400 ;
        RECT 0.2850 0.3075 0.3450 0.3675 ;
        RECT 0.1800 0.4800 0.2400 0.5400 ;
        RECT 0.0750 0.1725 0.1350 0.2325 ;
        RECT 0.0750 0.7875 0.1350 0.8475 ;
        LAYER M1 ;
        RECT 0.1575 0.1500 0.7950 0.2250 ;
        RECT 0.0525 0.1500 0.1575 0.2550 ;
    END
END OAI21_1010


MACRO OAI221_0011
    CLASS CORE ;
    FOREIGN OAI221_0011 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.5200 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 1.5600 0.8100 1.9200 0.8850 ;
        RECT 1.4850 0.7125 1.5600 0.8850 ;
        RECT 0.7725 0.7125 1.4850 0.7875 ;
        RECT 0.7725 0.2625 0.8025 0.4125 ;
        RECT 0.6975 0.2625 0.7725 0.9225 ;
        RECT 0.6675 0.7125 0.6975 0.9225 ;
        VIA 1.8075 0.8475 VIA12_square ;
        VIA 1.3650 0.7500 VIA12_square ;
        VIA 0.7500 0.3375 VIA12_square ;
        VIA 0.7200 0.8475 VIA12_square ;
        END
    END ZN
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.4025 0.5625 1.7175 0.6375 ;
        RECT 1.3275 0.4125 1.4025 0.6375 ;
        RECT 1.0125 0.4125 1.3275 0.4875 ;
        VIA 1.3650 0.5175 VIA12_square ;
        END
    END C
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 2.0325 0.4350 2.0625 0.5850 ;
        RECT 1.9575 0.2625 2.0325 0.5850 ;
        RECT 1.4925 0.2625 1.9575 0.3375 ;
        VIA 2.0100 0.5100 VIA12_square ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 2.2800 0.4125 2.4525 0.7350 ;
        RECT 1.7775 0.6600 2.2800 0.7350 ;
        RECT 1.7025 0.4650 1.7775 0.7350 ;
        RECT 1.6275 0.4650 1.7025 0.5700 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.8100 0.4725 0.9000 0.5625 ;
        RECT 0.7350 0.4725 0.8100 0.7350 ;
        RECT 0.2925 0.6600 0.7350 0.7350 ;
        RECT 0.2175 0.4950 0.2925 0.7350 ;
        RECT 0.1425 0.4950 0.2175 0.6825 ;
        RECT 0.0675 0.3675 0.1425 0.6825 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.5625 0.1125 1.0275 0.1875 ;
        RECT 0.5625 0.4500 0.5925 0.6000 ;
        RECT 0.4875 0.1125 0.5625 0.6000 ;
        VIA 0.5400 0.5250 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 2.2650 -0.0750 2.5200 0.0750 ;
        RECT 2.1450 -0.0750 2.2650 0.1875 ;
        RECT 1.8450 -0.0750 2.1450 0.0750 ;
        RECT 1.7250 -0.0750 1.8450 0.2250 ;
        RECT 0.0000 -0.0750 1.7250 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 2.4750 0.9750 2.5200 1.1250 ;
        RECT 2.3550 0.8100 2.4750 1.1250 ;
        RECT 1.6200 0.9750 2.3550 1.1250 ;
        RECT 1.5150 0.6750 1.6200 1.1250 ;
        RECT 1.2150 0.9750 1.5150 1.1250 ;
        RECT 1.0950 0.6675 1.2150 1.1250 ;
        RECT 1.0125 0.9750 1.0950 1.1250 ;
        RECT 0.9075 0.6375 1.0125 1.1250 ;
        RECT 0.1425 0.9750 0.9075 1.1250 ;
        RECT 0.0675 0.7875 0.1425 1.1250 ;
        RECT 0.0000 0.9750 0.0675 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 2.3850 0.2475 2.4450 0.3075 ;
        RECT 2.3850 0.8175 2.4450 0.8775 ;
        RECT 2.2800 0.4950 2.3400 0.5550 ;
        RECT 2.1750 0.1200 2.2350 0.1800 ;
        RECT 2.0700 0.4950 2.1300 0.5550 ;
        RECT 1.9650 0.2925 2.0250 0.3525 ;
        RECT 1.9650 0.8250 2.0250 0.8850 ;
        RECT 1.8600 0.4950 1.9200 0.5550 ;
        RECT 1.7550 0.1575 1.8150 0.2175 ;
        RECT 1.6500 0.4875 1.7100 0.5475 ;
        RECT 1.5450 0.3075 1.6050 0.3675 ;
        RECT 1.5450 0.7050 1.6050 0.7650 ;
        RECT 1.5450 0.8700 1.6050 0.9300 ;
        RECT 1.4400 0.4875 1.5000 0.5475 ;
        RECT 1.3350 0.1575 1.3950 0.2175 ;
        RECT 1.3350 0.7350 1.3950 0.7950 ;
        RECT 1.2300 0.4875 1.2900 0.5475 ;
        RECT 1.1250 0.3075 1.1850 0.3675 ;
        RECT 1.1250 0.6675 1.1850 0.7275 ;
        RECT 1.1250 0.8325 1.1850 0.8925 ;
        RECT 0.9150 0.1575 0.9750 0.2175 ;
        RECT 0.9150 0.6675 0.9750 0.7275 ;
        RECT 0.9150 0.8325 0.9750 0.8925 ;
        RECT 0.8100 0.4875 0.8700 0.5475 ;
        RECT 0.7050 0.3075 0.7650 0.3675 ;
        RECT 0.6000 0.4950 0.6600 0.5550 ;
        RECT 0.4950 0.1575 0.5550 0.2175 ;
        RECT 0.4950 0.8175 0.5550 0.8775 ;
        RECT 0.3900 0.4950 0.4500 0.5550 ;
        RECT 0.2850 0.3075 0.3450 0.3675 ;
        RECT 0.1800 0.4950 0.2400 0.5550 ;
        RECT 0.0750 0.1800 0.1350 0.2400 ;
        RECT 0.0750 0.8175 0.1350 0.8775 ;
        LAYER M1 ;
        RECT 2.3775 0.2175 2.4525 0.3375 ;
        RECT 2.0700 0.2625 2.3775 0.3375 ;
        RECT 1.8525 0.4575 2.1375 0.5850 ;
        RECT 1.7250 0.8100 2.0850 0.9000 ;
        RECT 1.9350 0.2625 2.0700 0.3750 ;
        RECT 1.0950 0.3000 1.9350 0.3750 ;
        RECT 1.2075 0.4650 1.5300 0.5700 ;
        RECT 1.2900 0.6675 1.4400 0.9000 ;
        RECT 0.1575 0.1500 1.4250 0.2250 ;
        RECT 0.2550 0.3000 0.9750 0.3825 ;
        RECT 0.4500 0.8100 0.8025 0.9000 ;
        RECT 0.3825 0.4650 0.6600 0.5850 ;
        RECT 0.0525 0.1500 0.1575 0.2625 ;
    END
END OAI221_0011


MACRO OAI221_0111
    CLASS CORE ;
    FOREIGN OAI221_0111 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.5200 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 1.8375 0.2850 2.1525 0.7275 ;
        VIA 1.9950 0.3450 VIA12_slot ;
        VIA 1.9950 0.6675 VIA12_slot ;
        END
    END ZN
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.6750 0.2625 1.1025 0.3375 ;
        RECT 0.6000 0.2625 0.6750 0.6375 ;
        RECT 0.5700 0.4875 0.6000 0.6375 ;
        VIA 0.6225 0.5625 VIA12_square ;
        END
    END C
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.7950 0.4125 1.2600 0.4875 ;
        VIA 1.1100 0.4500 VIA12_square ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.8250 0.5625 0.9825 0.6375 ;
        RECT 0.7500 0.5625 0.8250 0.9375 ;
        RECT 0.2850 0.8625 0.7500 0.9375 ;
        VIA 0.8700 0.6000 VIA12_square ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1575 0.4800 0.2625 0.5850 ;
        RECT 0.0525 0.3675 0.1575 0.6825 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.1650 0.7125 0.6300 0.7875 ;
        VIA 0.3600 0.7500 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 2.4525 -0.0750 2.5200 0.0750 ;
        RECT 2.3775 -0.0750 2.4525 0.3150 ;
        RECT 2.0550 -0.0750 2.3775 0.0750 ;
        RECT 1.9350 -0.0750 2.0550 0.1950 ;
        RECT 1.6350 -0.0750 1.9350 0.0750 ;
        RECT 1.5150 -0.0750 1.6350 0.1800 ;
        RECT 1.0050 -0.0750 1.5150 0.0750 ;
        RECT 0.8850 -0.0750 1.0050 0.1875 ;
        RECT 0.0000 -0.0750 0.8850 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 2.4525 0.9750 2.5200 1.1250 ;
        RECT 2.3775 0.6375 2.4525 1.1250 ;
        RECT 2.0325 0.9750 2.3775 1.1250 ;
        RECT 1.9575 0.8175 2.0325 1.1250 ;
        RECT 1.6350 0.9750 1.9575 1.1250 ;
        RECT 1.5150 0.8625 1.6350 1.1250 ;
        RECT 0.7950 0.9750 1.5150 1.1250 ;
        RECT 0.6750 0.8700 0.7950 1.1250 ;
        RECT 0.1650 0.9750 0.6750 1.1250 ;
        RECT 0.0450 0.8325 0.1650 1.1250 ;
        RECT 0.0000 0.9750 0.0450 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 2.3850 0.2250 2.4450 0.2850 ;
        RECT 2.3850 0.6675 2.4450 0.7275 ;
        RECT 2.3850 0.8325 2.4450 0.8925 ;
        RECT 2.2800 0.4650 2.3400 0.5250 ;
        RECT 2.1750 0.2250 2.2350 0.2850 ;
        RECT 2.1750 0.7200 2.2350 0.7800 ;
        RECT 2.0700 0.4650 2.1300 0.5250 ;
        RECT 1.9650 0.1275 2.0250 0.1875 ;
        RECT 1.9650 0.8475 2.0250 0.9075 ;
        RECT 1.8600 0.4650 1.9200 0.5250 ;
        RECT 1.7550 0.2250 1.8150 0.2850 ;
        RECT 1.7550 0.7200 1.8150 0.7800 ;
        RECT 1.6500 0.4650 1.7100 0.5250 ;
        RECT 1.5450 0.1200 1.6050 0.1800 ;
        RECT 1.5450 0.8625 1.6050 0.9225 ;
        RECT 1.4400 0.4650 1.5000 0.5250 ;
        RECT 1.3350 0.2175 1.3950 0.2775 ;
        RECT 1.3350 0.7650 1.3950 0.8250 ;
        RECT 1.1250 0.2325 1.1850 0.2925 ;
        RECT 1.1250 0.8175 1.1850 0.8775 ;
        RECT 1.0275 0.4800 1.0875 0.5400 ;
        RECT 0.9150 0.1275 0.9750 0.1875 ;
        RECT 0.8100 0.4800 0.8700 0.5400 ;
        RECT 0.7050 0.2325 0.7650 0.2925 ;
        RECT 0.7050 0.8700 0.7650 0.9300 ;
        RECT 0.6000 0.4950 0.6600 0.5550 ;
        RECT 0.4950 0.1650 0.5550 0.2250 ;
        RECT 0.4950 0.7500 0.5550 0.8100 ;
        RECT 0.3900 0.4950 0.4500 0.5550 ;
        RECT 0.2850 0.3225 0.3450 0.3825 ;
        RECT 0.1725 0.4950 0.2325 0.5550 ;
        RECT 0.0750 0.1950 0.1350 0.2550 ;
        RECT 0.0750 0.8325 0.1350 0.8925 ;
        LAYER M1 ;
        RECT 1.6725 0.4575 2.3700 0.5325 ;
        RECT 2.1525 0.1950 2.2575 0.3825 ;
        RECT 2.1675 0.6225 2.2425 0.8325 ;
        RECT 1.8225 0.6225 2.1675 0.7125 ;
        RECT 1.8375 0.2925 2.1525 0.3825 ;
        RECT 1.7475 0.1950 1.8375 0.3825 ;
        RECT 1.7475 0.6225 1.8225 0.8325 ;
        RECT 1.5975 0.2625 1.6725 0.7875 ;
        RECT 1.4175 0.2625 1.5975 0.3375 ;
        RECT 1.4175 0.7125 1.5975 0.7875 ;
        RECT 1.3125 0.4125 1.5225 0.6375 ;
        RECT 1.3125 0.1950 1.4175 0.3375 ;
        RECT 1.3125 0.7125 1.4175 0.8475 ;
        RECT 0.9450 0.7950 1.2075 0.9000 ;
        RECT 1.1100 0.1875 1.2000 0.3375 ;
        RECT 1.0275 0.4125 1.1925 0.6825 ;
        RECT 0.7800 0.2625 1.1100 0.3375 ;
        RECT 0.7875 0.4125 0.9525 0.6450 ;
        RECT 0.8700 0.7200 0.9450 0.9000 ;
        RECT 0.5625 0.7200 0.8700 0.7950 ;
        RECT 0.6900 0.1875 0.7800 0.3375 ;
        RECT 0.6075 0.4125 0.7125 0.6450 ;
        RECT 0.5550 0.4875 0.6075 0.6450 ;
        RECT 0.1575 0.1500 0.5850 0.2250 ;
        RECT 0.4875 0.7200 0.5625 0.8400 ;
        RECT 0.2325 0.3000 0.5325 0.4050 ;
        RECT 0.4125 0.4800 0.4800 0.5850 ;
        RECT 0.3375 0.4800 0.4125 0.8325 ;
        RECT 0.3075 0.6675 0.3375 0.8325 ;
        RECT 0.0525 0.1500 0.1575 0.2775 ;
        LAYER VIA1 ;
        RECT 1.4175 0.4725 1.4925 0.5475 ;
        RECT 1.0575 0.8175 1.1325 0.8925 ;
        RECT 0.4050 0.3150 0.4800 0.3900 ;
        LAYER M2 ;
        RECT 1.4175 0.1125 1.4925 0.8925 ;
        RECT 0.4950 0.1125 1.4175 0.1875 ;
        RECT 0.9825 0.8175 1.4175 0.8925 ;
        RECT 0.4200 0.1125 0.4950 0.4275 ;
        RECT 0.3900 0.2775 0.4200 0.4275 ;
    END
END OAI221_0111


MACRO OAI221_1000
    CLASS CORE ;
    FOREIGN OAI221_1000 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.4700 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 0.3825 0.5625 0.8475 0.6375 ;
        VIA 0.5925 0.6000 VIA12_square ;
        END
    END ZN
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.8475 0.1125 1.3125 0.1875 ;
        RECT 0.7725 0.1125 0.8475 0.4875 ;
        RECT 0.6375 0.4125 0.7725 0.4875 ;
        VIA 0.7575 0.4500 VIA12_square ;
        END
    END C
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.3275 0.4125 1.4025 0.6825 ;
        RECT 1.2225 0.4125 1.3275 0.5700 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.9675 0.4650 1.0425 0.9375 ;
        RECT 0.4425 0.8625 0.9675 0.9375 ;
        VIA 1.0050 0.5475 VIA12_square ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1575 0.4800 0.2325 0.6000 ;
        RECT 0.0525 0.3675 0.1575 0.6825 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.2475 0.7125 0.7125 0.7875 ;
        VIA 0.3600 0.7500 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.2150 -0.0750 1.4700 0.0750 ;
        RECT 1.0950 -0.0750 1.2150 0.1875 ;
        RECT 0.0000 -0.0750 1.0950 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.0050 0.9750 1.4700 1.1250 ;
        RECT 0.8850 0.8700 1.0050 1.1250 ;
        RECT 0.1650 0.9750 0.8850 1.1250 ;
        RECT 0.0450 0.8325 0.1650 1.1250 ;
        RECT 0.0000 0.9750 0.0450 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.3350 0.1575 1.3950 0.2175 ;
        RECT 1.3350 0.8175 1.3950 0.8775 ;
        RECT 1.2300 0.4800 1.2900 0.5400 ;
        RECT 1.1250 0.1275 1.1850 0.1875 ;
        RECT 1.0200 0.4800 1.0800 0.5400 ;
        RECT 0.9150 0.1800 0.9750 0.2400 ;
        RECT 0.9150 0.8700 0.9750 0.9300 ;
        RECT 0.8025 0.4950 0.8625 0.5550 ;
        RECT 0.7050 0.1575 0.7650 0.2175 ;
        RECT 0.7050 0.8175 0.7650 0.8775 ;
        RECT 0.4950 0.1575 0.5550 0.2175 ;
        RECT 0.4950 0.8175 0.5550 0.8775 ;
        RECT 0.3900 0.4950 0.4500 0.5550 ;
        RECT 0.2850 0.3075 0.3450 0.3675 ;
        RECT 0.1725 0.5100 0.2325 0.5700 ;
        RECT 0.0750 0.1950 0.1350 0.2550 ;
        RECT 0.0750 0.8325 0.1350 0.8925 ;
        LAYER M1 ;
        RECT 1.3050 0.1500 1.4250 0.3375 ;
        RECT 1.1550 0.7950 1.4175 0.9000 ;
        RECT 1.0050 0.2625 1.3050 0.3375 ;
        RECT 1.0800 0.7200 1.1550 0.9000 ;
        RECT 0.9375 0.4200 1.1475 0.6450 ;
        RECT 0.7950 0.7200 1.0800 0.7950 ;
        RECT 0.9000 0.1500 1.0050 0.3375 ;
        RECT 0.8250 0.4650 0.8625 0.6450 ;
        RECT 0.7050 0.3675 0.8250 0.6450 ;
        RECT 0.1575 0.1500 0.7950 0.2250 ;
        RECT 0.6300 0.7200 0.7950 0.9000 ;
        RECT 0.5550 0.3000 0.6300 0.9000 ;
        RECT 0.3675 0.3000 0.5550 0.3750 ;
        RECT 0.4725 0.7875 0.5550 0.9000 ;
        RECT 0.3975 0.4800 0.4800 0.5850 ;
        RECT 0.3075 0.4800 0.3975 0.8325 ;
        RECT 0.2475 0.3000 0.3675 0.4050 ;
        RECT 0.0525 0.1500 0.1575 0.2775 ;
    END
END OAI221_1000


MACRO OAI221_1010
    CLASS CORE ;
    FOREIGN OAI221_1010 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.4700 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 0.3825 0.5625 0.8475 0.6375 ;
        VIA 0.5925 0.6000 VIA12_square ;
        END
    END ZN
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.8475 0.1125 1.3125 0.1875 ;
        RECT 0.7725 0.1125 0.8475 0.4875 ;
        RECT 0.6375 0.4125 0.7725 0.4875 ;
        VIA 0.7575 0.4500 VIA12_square ;
        END
    END C
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.3275 0.4125 1.4025 0.6825 ;
        RECT 1.2225 0.4125 1.3275 0.5700 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.9675 0.4650 1.0425 0.9375 ;
        RECT 0.4425 0.8625 0.9675 0.9375 ;
        VIA 1.0050 0.5475 VIA12_square ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1575 0.4800 0.2625 0.5850 ;
        RECT 0.0525 0.3675 0.1575 0.6825 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.2475 0.7125 0.7125 0.7875 ;
        VIA 0.3600 0.7500 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.2150 -0.0750 1.4700 0.0750 ;
        RECT 1.0950 -0.0750 1.2150 0.1875 ;
        RECT 0.0000 -0.0750 1.0950 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.0050 0.9750 1.4700 1.1250 ;
        RECT 0.8850 0.8700 1.0050 1.1250 ;
        RECT 0.1650 0.9750 0.8850 1.1250 ;
        RECT 0.0450 0.8325 0.1650 1.1250 ;
        RECT 0.0000 0.9750 0.0450 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.3350 0.2325 1.3950 0.2925 ;
        RECT 1.3350 0.8175 1.3950 0.8775 ;
        RECT 1.2300 0.4800 1.2900 0.5400 ;
        RECT 1.1250 0.1275 1.1850 0.1875 ;
        RECT 1.0200 0.4800 1.0800 0.5400 ;
        RECT 0.9150 0.2325 0.9750 0.2925 ;
        RECT 0.9150 0.8700 0.9750 0.9300 ;
        RECT 0.8025 0.4950 0.8625 0.5550 ;
        RECT 0.7050 0.1650 0.7650 0.2250 ;
        RECT 0.7050 0.7275 0.7650 0.7875 ;
        RECT 0.4950 0.1650 0.5550 0.2250 ;
        RECT 0.4950 0.7275 0.5550 0.7875 ;
        RECT 0.3900 0.4950 0.4500 0.5550 ;
        RECT 0.2850 0.3225 0.3450 0.3825 ;
        RECT 0.1725 0.4950 0.2325 0.5550 ;
        RECT 0.0750 0.1950 0.1350 0.2550 ;
        RECT 0.0750 0.8325 0.1350 0.8925 ;
        LAYER M1 ;
        RECT 1.1550 0.7950 1.4175 0.9000 ;
        RECT 1.3200 0.1875 1.4100 0.3375 ;
        RECT 0.9900 0.2625 1.3200 0.3375 ;
        RECT 1.0800 0.7200 1.1550 0.9000 ;
        RECT 0.9375 0.4200 1.1475 0.6450 ;
        RECT 0.6300 0.7200 1.0800 0.7950 ;
        RECT 0.9000 0.1875 0.9900 0.3375 ;
        RECT 0.8100 0.4650 0.8625 0.6450 ;
        RECT 0.7050 0.3675 0.8100 0.6450 ;
        RECT 0.1575 0.1500 0.7950 0.2250 ;
        RECT 0.5625 0.3000 0.6300 0.7950 ;
        RECT 0.5550 0.3000 0.5625 0.8325 ;
        RECT 0.3675 0.3000 0.5550 0.3750 ;
        RECT 0.4875 0.6675 0.5550 0.8325 ;
        RECT 0.4125 0.4800 0.4800 0.5850 ;
        RECT 0.3375 0.4800 0.4125 0.8325 ;
        RECT 0.2625 0.3000 0.3675 0.4050 ;
        RECT 0.3075 0.6675 0.3375 0.8325 ;
        RECT 0.0525 0.1500 0.1575 0.2775 ;
    END
END OAI221_1010


MACRO OAI222_0011
    CLASS CORE ;
    FOREIGN OAI222_0011 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.9400 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 2.1525 0.7950 2.3025 0.9000 ;
        RECT 1.6200 0.8100 2.1525 0.8850 ;
        RECT 1.5450 0.7125 1.6200 0.8850 ;
        RECT 0.9750 0.7125 1.5450 0.7875 ;
        RECT 0.9000 0.3000 0.9750 0.8850 ;
        RECT 0.7800 0.3000 0.9000 0.3750 ;
        RECT 0.6375 0.7800 0.9000 0.8850 ;
        VIA 2.2275 0.8475 VIA12_square ;
        VIA 1.6950 0.8475 VIA12_square ;
        VIA 0.8925 0.3375 VIA12_square ;
        VIA 0.7200 0.8475 VIA12_square ;
        END
    END ZN
    PIN C2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 2.3625 0.4125 2.4675 0.6000 ;
        RECT 1.9125 0.4125 2.3625 0.4875 ;
        VIA 2.4150 0.5175 VIA12_square ;
        END
    END C2
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 2.7000 0.4125 2.8725 0.7350 ;
        RECT 2.1975 0.6600 2.7000 0.7350 ;
        RECT 2.1225 0.4650 2.1975 0.7350 ;
        RECT 2.0400 0.4650 2.1225 0.5700 ;
        END
    END C1
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.6725 0.5625 1.9950 0.6375 ;
        RECT 1.5975 0.4125 1.6725 0.6375 ;
        RECT 1.2825 0.4125 1.5975 0.4875 ;
        VIA 1.6350 0.5175 VIA12_square ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.1250 0.5625 1.4400 0.6375 ;
        RECT 1.0500 0.1125 1.1250 0.6375 ;
        RECT 0.7350 0.1125 1.0500 0.1875 ;
        VIA 1.0875 0.5175 VIA12_square ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.8100 0.4725 0.9000 0.5475 ;
        RECT 0.7350 0.4725 0.8100 0.7350 ;
        RECT 0.2925 0.6600 0.7350 0.7350 ;
        RECT 0.2175 0.4875 0.2925 0.7350 ;
        RECT 0.1425 0.4875 0.2175 0.6825 ;
        RECT 0.0675 0.3675 0.1425 0.6825 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.5400 0.1125 0.6150 0.5925 ;
        RECT 0.0750 0.1125 0.5400 0.1875 ;
        RECT 0.5100 0.4425 0.5400 0.5925 ;
        VIA 0.5625 0.5175 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 2.6850 -0.0750 2.9400 0.0750 ;
        RECT 2.5650 -0.0750 2.6850 0.1875 ;
        RECT 2.2650 -0.0750 2.5650 0.0750 ;
        RECT 2.1450 -0.0750 2.2650 0.2250 ;
        RECT 0.0000 -0.0750 2.1450 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 2.8950 0.9750 2.9400 1.1250 ;
        RECT 2.7750 0.8175 2.8950 1.1250 ;
        RECT 2.0325 0.9750 2.7750 1.1250 ;
        RECT 1.9575 0.6750 2.0325 1.1250 ;
        RECT 1.2150 0.9750 1.9575 1.1250 ;
        RECT 1.0950 0.6675 1.2150 1.1250 ;
        RECT 1.0125 0.9750 1.0950 1.1250 ;
        RECT 0.9075 0.6375 1.0125 1.1250 ;
        RECT 0.1425 0.9750 0.9075 1.1250 ;
        RECT 0.0675 0.7875 0.1425 1.1250 ;
        RECT 0.0000 0.9750 0.0675 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 2.8050 0.2325 2.8650 0.2925 ;
        RECT 2.8050 0.8175 2.8650 0.8775 ;
        RECT 2.7000 0.4950 2.7600 0.5550 ;
        RECT 2.5950 0.1200 2.6550 0.1800 ;
        RECT 2.4900 0.4950 2.5500 0.5550 ;
        RECT 2.3850 0.2925 2.4450 0.3525 ;
        RECT 2.3850 0.8250 2.4450 0.8850 ;
        RECT 2.2800 0.4950 2.3400 0.5550 ;
        RECT 2.1750 0.1575 2.2350 0.2175 ;
        RECT 2.0700 0.4875 2.1300 0.5475 ;
        RECT 1.9650 0.3075 2.0250 0.3675 ;
        RECT 1.9650 0.7050 2.0250 0.7650 ;
        RECT 1.9650 0.8700 2.0250 0.9300 ;
        RECT 1.8600 0.4875 1.9200 0.5475 ;
        RECT 1.7550 0.1575 1.8150 0.2175 ;
        RECT 1.6500 0.4950 1.7100 0.5550 ;
        RECT 1.5450 0.3075 1.6050 0.3675 ;
        RECT 1.5450 0.8250 1.6050 0.8850 ;
        RECT 1.4400 0.4950 1.5000 0.5550 ;
        RECT 1.3350 0.1575 1.3950 0.2175 ;
        RECT 1.2300 0.4875 1.2900 0.5475 ;
        RECT 1.1250 0.3075 1.1850 0.3675 ;
        RECT 1.1250 0.6675 1.1850 0.7275 ;
        RECT 1.1250 0.8325 1.1850 0.8925 ;
        RECT 0.9150 0.1575 0.9750 0.2175 ;
        RECT 0.9150 0.6675 0.9750 0.7275 ;
        RECT 0.9150 0.8325 0.9750 0.8925 ;
        RECT 0.8100 0.4800 0.8700 0.5400 ;
        RECT 0.7050 0.3075 0.7650 0.3675 ;
        RECT 0.6000 0.4950 0.6600 0.5550 ;
        RECT 0.4950 0.1575 0.5550 0.2175 ;
        RECT 0.4950 0.8250 0.5550 0.8850 ;
        RECT 0.3900 0.4950 0.4500 0.5550 ;
        RECT 0.2850 0.3075 0.3450 0.3675 ;
        RECT 0.1800 0.4950 0.2400 0.5550 ;
        RECT 0.0750 0.1800 0.1350 0.2400 ;
        RECT 0.0750 0.8175 0.1350 0.8775 ;
        LAYER M1 ;
        RECT 2.7975 0.2025 2.8725 0.3375 ;
        RECT 2.4825 0.2625 2.7975 0.3375 ;
        RECT 2.2725 0.4575 2.5575 0.5850 ;
        RECT 2.1450 0.8100 2.5125 0.9000 ;
        RECT 2.3475 0.2625 2.4825 0.3750 ;
        RECT 1.0950 0.3000 2.3475 0.3750 ;
        RECT 1.8675 0.4650 1.9500 0.5700 ;
        RECT 1.7925 0.4650 1.8675 0.7350 ;
        RECT 0.1575 0.1500 1.8450 0.2250 ;
        RECT 1.4100 0.8100 1.8075 0.9000 ;
        RECT 1.3650 0.6600 1.7925 0.7350 ;
        RECT 1.4400 0.4575 1.7100 0.5850 ;
        RECT 1.2900 0.4800 1.3650 0.7350 ;
        RECT 1.0050 0.4800 1.2900 0.5550 ;
        RECT 0.2550 0.3000 0.9750 0.3825 ;
        RECT 0.4500 0.8100 0.8025 0.9000 ;
        RECT 0.3825 0.4575 0.6600 0.5850 ;
        RECT 0.0525 0.1500 0.1575 0.2625 ;
    END
END OAI222_0011


MACRO OAI222_0111
    CLASS CORE ;
    FOREIGN OAI222_0111 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.7300 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 1.8375 0.2850 2.1525 0.7275 ;
        VIA 1.9950 0.3450 VIA12_slot ;
        VIA 1.9950 0.6675 VIA12_slot ;
        END
    END ZN
    PIN C2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.1550 0.5625 1.6200 0.6375 ;
        VIA 1.2675 0.6000 VIA12_square ;
        END
    END C2
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.2525 0.4125 1.7175 0.4875 ;
        VIA 1.5225 0.4500 VIA12_square ;
        END
    END C1
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.8850 0.1125 1.3500 0.1875 ;
        RECT 0.8100 0.1125 0.8850 0.6825 ;
        RECT 0.6525 0.5325 0.8100 0.6825 ;
        VIA 0.7050 0.6075 VIA12_square ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.0350 0.2625 1.5000 0.3375 ;
        RECT 0.9600 0.2625 1.0350 0.6600 ;
        VIA 0.9975 0.5475 VIA12_square ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1425 0.4800 0.2700 0.5850 ;
        RECT 0.0675 0.3675 0.1425 0.6825 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.4275 0.1125 0.6900 0.1875 ;
        RECT 0.3525 0.1125 0.4275 0.7125 ;
        RECT 0.1500 0.1125 0.3525 0.1875 ;
        VIA 0.3900 0.6000 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 2.4750 -0.0750 2.7300 0.0750 ;
        RECT 2.3700 -0.0750 2.4750 0.2175 ;
        RECT 2.0325 -0.0750 2.3700 0.0750 ;
        RECT 1.9275 -0.0750 2.0325 0.2175 ;
        RECT 1.6200 -0.0750 1.9275 0.0750 ;
        RECT 1.5225 -0.0750 1.6200 0.2325 ;
        RECT 1.2150 -0.0750 1.5225 0.0750 ;
        RECT 1.0950 -0.0750 1.2150 0.2550 ;
        RECT 0.0000 -0.0750 1.0950 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 2.4675 0.9750 2.7300 1.1250 ;
        RECT 2.3625 0.8175 2.4675 1.1250 ;
        RECT 2.0250 0.9750 2.3625 1.1250 ;
        RECT 1.9350 0.8175 2.0250 1.1250 ;
        RECT 1.6200 0.9750 1.9350 1.1250 ;
        RECT 1.5150 0.7950 1.6200 1.1250 ;
        RECT 1.0050 0.9750 1.5150 1.1250 ;
        RECT 0.8850 0.7575 1.0050 1.1250 ;
        RECT 0.1425 0.9750 0.8850 1.1250 ;
        RECT 0.0675 0.7875 0.1425 1.1250 ;
        RECT 0.0000 0.9750 0.0675 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 2.5950 0.2250 2.6550 0.2850 ;
        RECT 2.5950 0.8100 2.6550 0.8700 ;
        RECT 2.4825 0.4950 2.5425 0.5550 ;
        RECT 2.3850 0.1275 2.4450 0.1875 ;
        RECT 2.3850 0.8475 2.4450 0.9075 ;
        RECT 2.2725 0.4875 2.3325 0.5475 ;
        RECT 2.1750 0.1575 2.2350 0.2175 ;
        RECT 2.1750 0.7500 2.2350 0.8100 ;
        RECT 2.0700 0.4650 2.1300 0.5250 ;
        RECT 1.9650 0.1275 2.0250 0.1875 ;
        RECT 1.9650 0.8475 2.0250 0.9075 ;
        RECT 1.8600 0.4650 1.9200 0.5250 ;
        RECT 1.7550 0.2250 1.8150 0.2850 ;
        RECT 1.7550 0.7350 1.8150 0.7950 ;
        RECT 1.6500 0.4875 1.7100 0.5475 ;
        RECT 1.5450 0.1425 1.6050 0.2025 ;
        RECT 1.5450 0.8250 1.6050 0.8850 ;
        RECT 1.4400 0.4950 1.5000 0.5550 ;
        RECT 1.3350 0.2400 1.3950 0.3000 ;
        RECT 1.2300 0.4950 1.2900 0.5550 ;
        RECT 1.1250 0.1800 1.1850 0.2400 ;
        RECT 1.1250 0.8100 1.1850 0.8700 ;
        RECT 0.9150 0.1725 0.9750 0.2325 ;
        RECT 0.9150 0.7725 0.9750 0.8325 ;
        RECT 0.8175 0.5250 0.8775 0.5850 ;
        RECT 0.7050 0.3300 0.7650 0.3900 ;
        RECT 0.6000 0.5025 0.6600 0.5625 ;
        RECT 0.4950 0.1575 0.5550 0.2175 ;
        RECT 0.4950 0.8100 0.5550 0.8700 ;
        RECT 0.3900 0.4950 0.4500 0.5550 ;
        RECT 0.2850 0.3225 0.3450 0.3825 ;
        RECT 0.1800 0.4950 0.2400 0.5550 ;
        RECT 0.0750 0.1800 0.1350 0.2400 ;
        RECT 0.0750 0.8175 0.1350 0.8775 ;
        LAYER M1 ;
        RECT 2.6175 0.1950 2.6925 0.9000 ;
        RECT 2.5725 0.1950 2.6175 0.3750 ;
        RECT 2.5800 0.7800 2.6175 0.9000 ;
        RECT 2.3325 0.3000 2.5725 0.3750 ;
        RECT 2.4075 0.4500 2.5425 0.7125 ;
        RECT 2.2575 0.3000 2.3325 0.5775 ;
        RECT 2.1825 0.1500 2.2650 0.2250 ;
        RECT 2.2500 0.4575 2.2575 0.5775 ;
        RECT 2.1825 0.7275 2.2575 0.8325 ;
        RECT 1.7100 0.4575 2.2500 0.5325 ;
        RECT 2.1075 0.1500 2.1825 0.3825 ;
        RECT 2.1075 0.6225 2.1825 0.8325 ;
        RECT 1.8375 0.2925 2.1075 0.3825 ;
        RECT 1.8450 0.6225 2.1075 0.7125 ;
        RECT 1.7700 0.6225 1.8450 0.8325 ;
        RECT 1.7325 0.1950 1.8375 0.3825 ;
        RECT 1.7400 0.6975 1.7700 0.8325 ;
        RECT 1.6350 0.4575 1.7100 0.5775 ;
        RECT 1.4850 0.3375 1.5600 0.7200 ;
        RECT 1.4100 0.4800 1.4850 0.7200 ;
        RECT 1.3200 0.2100 1.4100 0.4050 ;
        RECT 1.0950 0.7950 1.3950 0.9000 ;
        RECT 0.9300 0.3300 1.3200 0.4050 ;
        RECT 1.1700 0.4800 1.3200 0.7200 ;
        RECT 0.9225 0.4950 1.0950 0.6000 ;
        RECT 0.8925 0.1500 0.9975 0.2550 ;
        RECT 0.8100 0.3300 0.9300 0.4200 ;
        RECT 0.8175 0.4950 0.9225 0.6225 ;
        RECT 0.1575 0.1500 0.8925 0.2250 ;
        RECT 0.7050 0.3000 0.8100 0.4200 ;
        RECT 0.4500 0.8100 0.7800 0.9000 ;
        RECT 0.5625 0.4950 0.7425 0.7125 ;
        RECT 0.2625 0.3000 0.6300 0.4050 ;
        RECT 0.3450 0.4800 0.4875 0.7350 ;
        RECT 0.0525 0.1500 0.1575 0.2625 ;
        LAYER VIA1 ;
        RECT 2.4075 0.5625 2.4825 0.6375 ;
        RECT 1.1850 0.8100 1.2600 0.8850 ;
        RECT 0.6450 0.8100 0.7200 0.8850 ;
        RECT 0.5025 0.3150 0.5775 0.3900 ;
        LAYER M2 ;
        RECT 2.3775 0.5625 2.5575 0.6375 ;
        RECT 2.3025 0.5625 2.3775 0.9375 ;
        RECT 1.3575 0.8625 2.3025 0.9375 ;
        RECT 1.2825 0.8100 1.3575 0.9375 ;
        RECT 0.5775 0.8100 1.2825 0.8850 ;
        RECT 0.5775 0.2700 0.6075 0.3750 ;
        RECT 0.5025 0.2700 0.5775 0.8850 ;
    END
END OAI222_0111


MACRO OAI222_1000
    CLASS CORE ;
    FOREIGN OAI222_1000 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.6800 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 0.8625 0.7125 1.0125 0.8775 ;
        RECT 0.3975 0.7125 0.8625 0.7875 ;
        VIA 0.9375 0.8250 VIA12_square ;
        VIA 0.5625 0.7500 VIA12_square ;
        END
    END ZN
    PIN C2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.1325 0.7125 1.5975 0.7875 ;
        VIA 1.3350 0.7500 VIA12_square ;
        END
    END C2
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.5225 0.4125 1.6275 0.6825 ;
        RECT 1.4475 0.4125 1.5225 0.5850 ;
        END
    END C1
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.0500 0.1125 1.5150 0.1875 ;
        RECT 1.0500 0.4500 1.1400 0.5550 ;
        RECT 0.9750 0.1125 1.0500 0.5550 ;
        VIA 1.0575 0.5025 VIA12_square ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.8175 0.1125 0.8925 0.5700 ;
        RECT 0.3525 0.1125 0.8175 0.1875 ;
        RECT 0.7275 0.4650 0.8175 0.5700 ;
        VIA 0.8100 0.5175 VIA12_square ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1425 0.4575 0.2325 0.6825 ;
        RECT 0.0675 0.3675 0.1425 0.6825 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.4650 0.2625 0.6975 0.3375 ;
        RECT 0.3600 0.2625 0.4650 0.6150 ;
        RECT 0.1125 0.2625 0.3600 0.3375 ;
        VIA 0.4125 0.5325 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.4250 -0.0750 1.6800 0.0750 ;
        RECT 1.3050 -0.0750 1.4250 0.1875 ;
        RECT 0.0000 -0.0750 1.3050 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.6125 0.9750 1.6800 1.1250 ;
        RECT 1.5075 0.8025 1.6125 1.1250 ;
        RECT 0.7875 0.9750 1.5075 1.1250 ;
        RECT 0.6825 0.8025 0.7875 1.1250 ;
        RECT 0.1425 0.9750 0.6825 1.1250 ;
        RECT 0.0675 0.7875 0.1425 1.1250 ;
        RECT 0.0000 0.9750 0.0675 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.5450 0.1575 1.6050 0.2175 ;
        RECT 1.5450 0.8325 1.6050 0.8925 ;
        RECT 1.4475 0.4800 1.5075 0.5400 ;
        RECT 1.3350 0.1200 1.3950 0.1800 ;
        RECT 1.2375 0.4950 1.2975 0.5550 ;
        RECT 1.1250 0.1800 1.1850 0.2400 ;
        RECT 1.1250 0.8100 1.1850 0.8700 ;
        RECT 1.0200 0.4950 1.0800 0.5550 ;
        RECT 0.9150 0.1575 0.9750 0.2175 ;
        RECT 0.8100 0.4950 0.8700 0.5550 ;
        RECT 0.7050 0.3075 0.7650 0.3675 ;
        RECT 0.7050 0.8325 0.7650 0.8925 ;
        RECT 0.4950 0.1575 0.5550 0.2175 ;
        RECT 0.4950 0.8250 0.5550 0.8850 ;
        RECT 0.3900 0.4950 0.4500 0.5550 ;
        RECT 0.2850 0.3075 0.3450 0.3675 ;
        RECT 0.1725 0.4950 0.2325 0.5550 ;
        RECT 0.0750 0.1725 0.1350 0.2325 ;
        RECT 0.0750 0.8175 0.1350 0.8775 ;
        LAYER M1 ;
        RECT 1.5150 0.1500 1.6350 0.3375 ;
        RECT 1.2150 0.2625 1.5150 0.3375 ;
        RECT 1.3725 0.6675 1.4025 0.8325 ;
        RECT 1.2900 0.4575 1.3725 0.8325 ;
        RECT 1.2375 0.4575 1.2900 0.5925 ;
        RECT 1.1925 0.1500 1.2150 0.3375 ;
        RECT 0.8625 0.7725 1.2150 0.9000 ;
        RECT 1.1100 0.1500 1.1925 0.3750 ;
        RECT 0.9750 0.4500 1.1625 0.6825 ;
        RECT 0.7875 0.3000 1.1100 0.3750 ;
        RECT 0.1575 0.1500 1.0050 0.2250 ;
        RECT 0.6825 0.4800 0.9000 0.6825 ;
        RECT 0.6750 0.3000 0.7875 0.4050 ;
        RECT 0.5250 0.3000 0.6000 0.9000 ;
        RECT 0.2550 0.3000 0.5250 0.3750 ;
        RECT 0.4275 0.7875 0.5250 0.9000 ;
        RECT 0.3075 0.4500 0.4500 0.7125 ;
        RECT 0.0525 0.1500 0.1575 0.2550 ;
    END
END OAI222_1000


MACRO OAI222_1010
    CLASS CORE ;
    FOREIGN OAI222_1010 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.6800 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 0.8625 0.7125 1.0125 0.8775 ;
        RECT 0.3975 0.7125 0.8625 0.7875 ;
        VIA 0.9375 0.8250 VIA12_square ;
        VIA 0.5625 0.7500 VIA12_square ;
        END
    END ZN
    PIN C2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.1325 0.7125 1.5975 0.7875 ;
        VIA 1.3350 0.7500 VIA12_square ;
        END
    END C2
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.5225 0.4125 1.6275 0.6825 ;
        RECT 1.4475 0.4125 1.5225 0.5850 ;
        END
    END C1
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.0500 0.1125 1.5150 0.1875 ;
        RECT 1.0500 0.4500 1.1400 0.5550 ;
        RECT 0.9750 0.1125 1.0500 0.5550 ;
        VIA 1.0575 0.5025 VIA12_square ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.8175 0.1125 0.8925 0.5700 ;
        RECT 0.3525 0.1125 0.8175 0.1875 ;
        RECT 0.7275 0.4650 0.8175 0.5700 ;
        VIA 0.8100 0.5175 VIA12_square ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1425 0.4575 0.2325 0.6825 ;
        RECT 0.0675 0.3675 0.1425 0.6825 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.4650 0.2625 0.6975 0.3375 ;
        RECT 0.3600 0.2625 0.4650 0.6150 ;
        RECT 0.1125 0.2625 0.3600 0.3375 ;
        VIA 0.4125 0.5325 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.4250 -0.0750 1.6800 0.0750 ;
        RECT 1.3050 -0.0750 1.4250 0.1875 ;
        RECT 0.0000 -0.0750 1.3050 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.6125 0.9750 1.6800 1.1250 ;
        RECT 1.5075 0.8025 1.6125 1.1250 ;
        RECT 0.7875 0.9750 1.5075 1.1250 ;
        RECT 0.6825 0.8025 0.7875 1.1250 ;
        RECT 0.1425 0.9750 0.6825 1.1250 ;
        RECT 0.0675 0.7875 0.1425 1.1250 ;
        RECT 0.0000 0.9750 0.0675 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.5450 0.1575 1.6050 0.2175 ;
        RECT 1.5450 0.8325 1.6050 0.8925 ;
        RECT 1.4475 0.4800 1.5075 0.5400 ;
        RECT 1.3350 0.1200 1.3950 0.1800 ;
        RECT 1.2375 0.4950 1.2975 0.5550 ;
        RECT 1.1250 0.1800 1.1850 0.2400 ;
        RECT 1.1250 0.8100 1.1850 0.8700 ;
        RECT 1.0200 0.4950 1.0800 0.5550 ;
        RECT 0.9150 0.1575 0.9750 0.2175 ;
        RECT 0.8100 0.4950 0.8700 0.5550 ;
        RECT 0.7050 0.3075 0.7650 0.3675 ;
        RECT 0.7050 0.8325 0.7650 0.8925 ;
        RECT 0.4950 0.1575 0.5550 0.2175 ;
        RECT 0.4950 0.8250 0.5550 0.8850 ;
        RECT 0.3900 0.4950 0.4500 0.5550 ;
        RECT 0.2850 0.3075 0.3450 0.3675 ;
        RECT 0.1725 0.4950 0.2325 0.5550 ;
        RECT 0.0750 0.1725 0.1350 0.2325 ;
        RECT 0.0750 0.8175 0.1350 0.8775 ;
        LAYER M1 ;
        RECT 1.5150 0.1500 1.6350 0.3375 ;
        RECT 1.2150 0.2625 1.5150 0.3375 ;
        RECT 1.3725 0.6675 1.4025 0.8325 ;
        RECT 1.2900 0.4575 1.3725 0.8325 ;
        RECT 1.2375 0.4575 1.2900 0.5925 ;
        RECT 1.1925 0.1500 1.2150 0.3375 ;
        RECT 0.8625 0.7725 1.2150 0.9000 ;
        RECT 1.1100 0.1500 1.1925 0.3750 ;
        RECT 0.9750 0.4500 1.1625 0.6825 ;
        RECT 0.7875 0.3000 1.1100 0.3750 ;
        RECT 0.1575 0.1500 1.0050 0.2250 ;
        RECT 0.6825 0.4800 0.9000 0.6825 ;
        RECT 0.6750 0.3000 0.7875 0.4050 ;
        RECT 0.5250 0.3000 0.6000 0.9000 ;
        RECT 0.2550 0.3000 0.5250 0.3750 ;
        RECT 0.4275 0.7875 0.5250 0.9000 ;
        RECT 0.3075 0.4500 0.4500 0.7125 ;
        RECT 0.0525 0.1500 0.1575 0.2550 ;
    END
END OAI222_1010


MACRO OAI22_0011
    CLASS CORE ;
    FOREIGN OAI22_0011 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.6100 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 1.1025 0.6525 3.9375 0.7725 ;
        RECT 1.1025 0.2775 1.2600 0.3975 ;
        RECT 0.7875 0.2775 1.1025 0.7725 ;
        RECT 0.6300 0.2775 0.7875 0.3975 ;
        RECT 0.6300 0.6525 0.7875 0.7725 ;
        VIA 3.7800 0.7125 VIA12_slot ;
        VIA 1.1025 0.7125 VIA12_slot ;
        VIA 1.1025 0.3375 VIA12_slot ;
        VIA 0.7875 0.3375 VIA12_slot ;
        VIA 0.7875 0.7125 VIA12_slot ;
        END
    END ZN
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 8.3100 0.4125 8.4750 0.6375 ;
        RECT 6.0375 0.4725 8.3100 0.5775 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 5.7675 0.4125 5.9325 0.6375 ;
        RECT 3.5100 0.4575 5.7675 0.5625 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 3.4050 0.4125 3.7575 0.4875 ;
        RECT 3.2700 0.4125 3.4050 0.5775 ;
        VIA 3.3375 0.5025 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1425 0.4950 1.7325 0.5850 ;
        RECT 0.0375 0.3675 0.1425 0.6825 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 8.3550 -0.0750 8.6100 0.0750 ;
        RECT 8.2350 -0.0750 8.3550 0.1875 ;
        RECT 7.9350 -0.0750 8.2350 0.0750 ;
        RECT 7.8150 -0.0750 7.9350 0.1875 ;
        RECT 7.5150 -0.0750 7.8150 0.0750 ;
        RECT 7.3950 -0.0750 7.5150 0.1875 ;
        RECT 7.0950 -0.0750 7.3950 0.0750 ;
        RECT 6.9750 -0.0750 7.0950 0.1875 ;
        RECT 6.6750 -0.0750 6.9750 0.0750 ;
        RECT 6.5550 -0.0750 6.6750 0.1875 ;
        RECT 6.2550 -0.0750 6.5550 0.0750 ;
        RECT 6.1350 -0.0750 6.2550 0.1875 ;
        RECT 5.8350 -0.0750 6.1350 0.0750 ;
        RECT 5.7150 -0.0750 5.8350 0.1875 ;
        RECT 5.4150 -0.0750 5.7150 0.0750 ;
        RECT 5.2950 -0.0750 5.4150 0.1875 ;
        RECT 4.9950 -0.0750 5.2950 0.0750 ;
        RECT 4.8750 -0.0750 4.9950 0.1875 ;
        RECT 4.5750 -0.0750 4.8750 0.0750 ;
        RECT 4.4550 -0.0750 4.5750 0.1875 ;
        RECT 4.1550 -0.0750 4.4550 0.0750 ;
        RECT 4.0350 -0.0750 4.1550 0.1875 ;
        RECT 3.7500 -0.0750 4.0350 0.0750 ;
        RECT 3.6150 -0.0750 3.7500 0.1875 ;
        RECT 0.0000 -0.0750 3.6150 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 8.3550 0.9750 8.6100 1.1250 ;
        RECT 8.2350 0.8625 8.3550 1.1250 ;
        RECT 7.9350 0.9750 8.2350 1.1250 ;
        RECT 7.8150 0.8625 7.9350 1.1250 ;
        RECT 7.5150 0.9750 7.8150 1.1250 ;
        RECT 7.3950 0.8625 7.5150 1.1250 ;
        RECT 7.0950 0.9750 7.3950 1.1250 ;
        RECT 6.9750 0.8625 7.0950 1.1250 ;
        RECT 6.6750 0.9750 6.9750 1.1250 ;
        RECT 6.5550 0.8625 6.6750 1.1250 ;
        RECT 6.2550 0.9750 6.5550 1.1250 ;
        RECT 6.1350 0.8625 6.2550 1.1250 ;
        RECT 3.3150 0.9750 6.1350 1.1250 ;
        RECT 3.1950 0.8250 3.3150 1.1250 ;
        RECT 2.8950 0.9750 3.1950 1.1250 ;
        RECT 2.7750 0.8250 2.8950 1.1250 ;
        RECT 2.4750 0.9750 2.7750 1.1250 ;
        RECT 2.3550 0.8250 2.4750 1.1250 ;
        RECT 2.0550 0.9750 2.3550 1.1250 ;
        RECT 1.9350 0.8250 2.0550 1.1250 ;
        RECT 0.0000 0.9750 1.9350 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 8.4750 0.2325 8.5350 0.2925 ;
        RECT 8.4750 0.7575 8.5350 0.8175 ;
        RECT 8.3700 0.4950 8.4300 0.5550 ;
        RECT 8.2650 0.1275 8.3250 0.1875 ;
        RECT 8.2650 0.8625 8.3250 0.9225 ;
        RECT 8.1600 0.4950 8.2200 0.5550 ;
        RECT 8.0550 0.2700 8.1150 0.3300 ;
        RECT 8.0550 0.7200 8.1150 0.7800 ;
        RECT 7.9500 0.4950 8.0100 0.5550 ;
        RECT 7.8450 0.1275 7.9050 0.1875 ;
        RECT 7.8450 0.8625 7.9050 0.9225 ;
        RECT 7.7400 0.4950 7.8000 0.5550 ;
        RECT 7.6350 0.2700 7.6950 0.3300 ;
        RECT 7.6350 0.7200 7.6950 0.7800 ;
        RECT 7.5300 0.4950 7.5900 0.5550 ;
        RECT 7.4250 0.1275 7.4850 0.1875 ;
        RECT 7.4250 0.8625 7.4850 0.9225 ;
        RECT 7.3200 0.4950 7.3800 0.5550 ;
        RECT 7.2150 0.2700 7.2750 0.3300 ;
        RECT 7.2150 0.7200 7.2750 0.7800 ;
        RECT 7.1100 0.4950 7.1700 0.5550 ;
        RECT 7.0050 0.1275 7.0650 0.1875 ;
        RECT 7.0050 0.8625 7.0650 0.9225 ;
        RECT 6.9000 0.4950 6.9600 0.5550 ;
        RECT 6.7950 0.2700 6.8550 0.3300 ;
        RECT 6.7950 0.7200 6.8550 0.7800 ;
        RECT 6.6900 0.4950 6.7500 0.5550 ;
        RECT 6.5850 0.1275 6.6450 0.1875 ;
        RECT 6.5850 0.8625 6.6450 0.9225 ;
        RECT 6.4800 0.4950 6.5400 0.5550 ;
        RECT 6.3750 0.2700 6.4350 0.3300 ;
        RECT 6.3750 0.7200 6.4350 0.7800 ;
        RECT 6.2700 0.4950 6.3300 0.5550 ;
        RECT 6.1650 0.1275 6.2250 0.1875 ;
        RECT 6.1650 0.8625 6.2250 0.9225 ;
        RECT 6.0600 0.4950 6.1200 0.5550 ;
        RECT 5.9550 0.2700 6.0150 0.3300 ;
        RECT 5.9550 0.7725 6.0150 0.8325 ;
        RECT 5.8500 0.5100 5.9100 0.5700 ;
        RECT 5.7450 0.1275 5.8050 0.1875 ;
        RECT 5.6400 0.4800 5.7000 0.5400 ;
        RECT 5.5350 0.2700 5.5950 0.3300 ;
        RECT 5.5350 0.6900 5.5950 0.7500 ;
        RECT 5.4300 0.4800 5.4900 0.5400 ;
        RECT 5.3250 0.1275 5.3850 0.1875 ;
        RECT 5.3250 0.8325 5.3850 0.8925 ;
        RECT 5.2200 0.4800 5.2800 0.5400 ;
        RECT 5.1150 0.2700 5.1750 0.3300 ;
        RECT 5.1150 0.6900 5.1750 0.7500 ;
        RECT 5.0100 0.4800 5.0700 0.5400 ;
        RECT 4.9050 0.1275 4.9650 0.1875 ;
        RECT 4.9050 0.8325 4.9650 0.8925 ;
        RECT 4.8000 0.4800 4.8600 0.5400 ;
        RECT 4.6950 0.2700 4.7550 0.3300 ;
        RECT 4.6950 0.6900 4.7550 0.7500 ;
        RECT 4.5900 0.4800 4.6500 0.5400 ;
        RECT 4.4850 0.1275 4.5450 0.1875 ;
        RECT 4.4850 0.8325 4.5450 0.8925 ;
        RECT 4.3800 0.4800 4.4400 0.5400 ;
        RECT 4.2750 0.2700 4.3350 0.3300 ;
        RECT 4.2750 0.6900 4.3350 0.7500 ;
        RECT 4.1700 0.4800 4.2300 0.5400 ;
        RECT 4.0650 0.1275 4.1250 0.1875 ;
        RECT 4.0650 0.8325 4.1250 0.8925 ;
        RECT 3.9600 0.4800 4.0200 0.5400 ;
        RECT 3.8550 0.2700 3.9150 0.3300 ;
        RECT 3.8550 0.6900 3.9150 0.7500 ;
        RECT 3.7500 0.4800 3.8100 0.5400 ;
        RECT 3.6450 0.1275 3.7050 0.1875 ;
        RECT 3.5400 0.4725 3.6000 0.5325 ;
        RECT 3.4350 0.2100 3.4950 0.2700 ;
        RECT 3.4350 0.7575 3.4950 0.8175 ;
        RECT 3.3300 0.5100 3.3900 0.5700 ;
        RECT 3.2250 0.3075 3.2850 0.3675 ;
        RECT 3.2250 0.8400 3.2850 0.9000 ;
        RECT 3.1200 0.5100 3.1800 0.5700 ;
        RECT 3.0150 0.1575 3.0750 0.2175 ;
        RECT 3.0150 0.7575 3.0750 0.8175 ;
        RECT 2.9100 0.5100 2.9700 0.5700 ;
        RECT 2.8050 0.3075 2.8650 0.3675 ;
        RECT 2.8050 0.8400 2.8650 0.9000 ;
        RECT 2.7000 0.5100 2.7600 0.5700 ;
        RECT 2.5950 0.1575 2.6550 0.2175 ;
        RECT 2.5950 0.7575 2.6550 0.8175 ;
        RECT 2.4900 0.5100 2.5500 0.5700 ;
        RECT 2.3850 0.3075 2.4450 0.3675 ;
        RECT 2.3850 0.8400 2.4450 0.9000 ;
        RECT 2.2800 0.5100 2.3400 0.5700 ;
        RECT 2.1750 0.1575 2.2350 0.2175 ;
        RECT 2.1750 0.7575 2.2350 0.8175 ;
        RECT 2.0700 0.5100 2.1300 0.5700 ;
        RECT 1.9650 0.3075 2.0250 0.3675 ;
        RECT 1.9650 0.8400 2.0250 0.9000 ;
        RECT 1.8675 0.5100 1.9275 0.5700 ;
        RECT 1.7550 0.1575 1.8150 0.2175 ;
        RECT 1.7550 0.7650 1.8150 0.8250 ;
        RECT 1.6425 0.5025 1.7025 0.5625 ;
        RECT 1.5450 0.3075 1.6050 0.3675 ;
        RECT 1.5450 0.6825 1.6050 0.7425 ;
        RECT 1.4400 0.5025 1.5000 0.5625 ;
        RECT 1.3350 0.1650 1.3950 0.2250 ;
        RECT 1.3350 0.8325 1.3950 0.8925 ;
        RECT 1.2300 0.5025 1.2900 0.5625 ;
        RECT 1.1250 0.3075 1.1850 0.3675 ;
        RECT 1.1250 0.6825 1.1850 0.7425 ;
        RECT 1.0200 0.5025 1.0800 0.5625 ;
        RECT 0.9150 0.1650 0.9750 0.2250 ;
        RECT 0.9150 0.8325 0.9750 0.8925 ;
        RECT 0.8100 0.5025 0.8700 0.5625 ;
        RECT 0.7050 0.3075 0.7650 0.3675 ;
        RECT 0.7050 0.6825 0.7650 0.7425 ;
        RECT 0.6000 0.5100 0.6600 0.5700 ;
        RECT 0.4950 0.1650 0.5550 0.2250 ;
        RECT 0.4950 0.8325 0.5550 0.8925 ;
        RECT 0.3900 0.5100 0.4500 0.5700 ;
        RECT 0.2850 0.3225 0.3450 0.3825 ;
        RECT 0.2850 0.6825 0.3450 0.7425 ;
        RECT 0.1800 0.5100 0.2400 0.5700 ;
        RECT 0.0750 0.1725 0.1350 0.2325 ;
        RECT 0.0750 0.8175 0.1350 0.8775 ;
        LAYER M1 ;
        RECT 8.4675 0.1875 8.5425 0.3375 ;
        RECT 8.4675 0.7125 8.5425 0.8625 ;
        RECT 3.5025 0.2625 8.4675 0.3375 ;
        RECT 6.0225 0.7125 8.4675 0.7875 ;
        RECT 5.9475 0.7125 6.0225 0.9000 ;
        RECT 4.0200 0.8250 5.9475 0.9000 ;
        RECT 3.6075 0.6750 5.6400 0.7500 ;
        RECT 3.4275 0.1500 3.5025 0.3375 ;
        RECT 3.4275 0.6750 3.5025 0.8625 ;
        RECT 0.1575 0.1500 3.4275 0.2250 ;
        RECT 3.0825 0.6750 3.4275 0.7500 ;
        RECT 3.2550 0.4500 3.4200 0.5775 ;
        RECT 0.3825 0.3000 3.3150 0.3750 ;
        RECT 1.8375 0.5025 3.2550 0.5775 ;
        RECT 3.0075 0.6750 3.0825 0.8625 ;
        RECT 2.6625 0.6750 3.0075 0.7500 ;
        RECT 2.5875 0.6750 2.6625 0.8625 ;
        RECT 2.2425 0.6750 2.5875 0.7500 ;
        RECT 2.1675 0.6750 2.2425 0.8625 ;
        RECT 1.8225 0.6750 2.1675 0.7500 ;
        RECT 1.7475 0.6750 1.8225 0.9000 ;
        RECT 0.1575 0.8250 1.7475 0.9000 ;
        RECT 0.2550 0.6600 1.6425 0.7500 ;
        RECT 0.2625 0.3000 0.3825 0.4050 ;
        RECT 0.0525 0.1500 0.1575 0.2550 ;
        RECT 0.0525 0.7950 0.1575 0.9000 ;
        LAYER M2 ;
        RECT 1.1325 0.6525 3.9375 0.7725 ;
        RECT 1.1325 0.2775 1.2600 0.3975 ;
        RECT 0.6300 0.2775 0.7575 0.3975 ;
        RECT 0.6300 0.6525 0.7575 0.7725 ;
    END
END OAI22_0011


MACRO OAI22_0111
    CLASS CORE ;
    FOREIGN OAI22_0111 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.7800 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 0.3675 0.2925 0.6825 0.7725 ;
        VIA 0.5250 0.3525 VIA12_slot ;
        VIA 0.5250 0.7125 VIA12_slot ;
        END
    END ZN
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 3.6075 0.3675 3.7125 0.6375 ;
        RECT 3.5475 0.4725 3.6075 0.6375 ;
        RECT 2.8800 0.4725 3.5475 0.5775 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 2.6625 0.4125 2.9775 0.4875 ;
        RECT 2.5875 0.4125 2.6625 0.6375 ;
        RECT 2.2725 0.5625 2.5875 0.6375 ;
        VIA 2.6250 0.5250 VIA12_square ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.4625 0.5625 1.7775 0.6375 ;
        RECT 1.3875 0.4125 1.4625 0.6375 ;
        RECT 1.0725 0.4125 1.3875 0.4875 ;
        VIA 1.4250 0.5250 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.9225 0.7125 1.3875 0.7875 ;
        RECT 0.8475 0.4500 0.9225 0.7875 ;
        RECT 0.7875 0.4500 0.8475 0.6000 ;
        VIA 0.8400 0.5250 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 3.7275 -0.0750 3.7800 0.0750 ;
        RECT 3.6225 -0.0750 3.7275 0.2400 ;
        RECT 3.3150 -0.0750 3.6225 0.0750 ;
        RECT 3.1950 -0.0750 3.3150 0.2400 ;
        RECT 2.8950 -0.0750 3.1950 0.0750 ;
        RECT 2.7750 -0.0750 2.8950 0.2400 ;
        RECT 2.4750 -0.0750 2.7750 0.0750 ;
        RECT 2.3550 -0.0750 2.4750 0.2400 ;
        RECT 2.0400 -0.0750 2.3550 0.0750 ;
        RECT 1.9500 -0.0750 2.0400 0.3150 ;
        RECT 0.0000 -0.0750 1.9500 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 3.5250 0.9750 3.7800 1.1250 ;
        RECT 3.4050 0.8625 3.5250 1.1250 ;
        RECT 3.0975 0.9750 3.4050 1.1250 ;
        RECT 2.9925 0.8100 3.0975 1.1250 ;
        RECT 1.6275 0.9750 2.9925 1.1250 ;
        RECT 1.5225 0.8250 1.6275 1.1250 ;
        RECT 1.2075 0.9750 1.5225 1.1250 ;
        RECT 1.1025 0.8250 1.2075 1.1250 ;
        RECT 0.0000 0.9750 1.1025 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 3.6450 0.1575 3.7050 0.2175 ;
        RECT 3.6450 0.7575 3.7050 0.8175 ;
        RECT 3.5400 0.4950 3.6000 0.5550 ;
        RECT 3.4350 0.2400 3.4950 0.3000 ;
        RECT 3.4350 0.8700 3.4950 0.9300 ;
        RECT 3.3300 0.4950 3.3900 0.5550 ;
        RECT 3.2250 0.1725 3.2850 0.2325 ;
        RECT 3.2250 0.6975 3.2850 0.7575 ;
        RECT 3.1200 0.4950 3.1800 0.5550 ;
        RECT 3.0150 0.2400 3.0750 0.3000 ;
        RECT 3.0150 0.8325 3.0750 0.8925 ;
        RECT 2.9100 0.4950 2.9700 0.5550 ;
        RECT 2.8050 0.1725 2.8650 0.2325 ;
        RECT 2.8050 0.7575 2.8650 0.8175 ;
        RECT 2.7000 0.4950 2.7600 0.5550 ;
        RECT 2.5950 0.2400 2.6550 0.3000 ;
        RECT 2.5950 0.8175 2.6550 0.8775 ;
        RECT 2.4900 0.4950 2.5500 0.5550 ;
        RECT 2.3850 0.1725 2.4450 0.2325 ;
        RECT 2.3850 0.6750 2.4450 0.7350 ;
        RECT 2.2800 0.4950 2.3400 0.5550 ;
        RECT 2.1750 0.2400 2.2350 0.3000 ;
        RECT 2.1750 0.8175 2.2350 0.8775 ;
        RECT 2.0700 0.4950 2.1300 0.5550 ;
        RECT 1.9650 0.2175 2.0250 0.2775 ;
        RECT 1.9650 0.7575 2.0250 0.8175 ;
        RECT 1.7550 0.2550 1.8150 0.3150 ;
        RECT 1.7550 0.7575 1.8150 0.8175 ;
        RECT 1.6500 0.4950 1.7100 0.5550 ;
        RECT 1.5450 0.1725 1.6050 0.2325 ;
        RECT 1.5450 0.8475 1.6050 0.9075 ;
        RECT 1.4400 0.4950 1.5000 0.5550 ;
        RECT 1.3350 0.3225 1.3950 0.3825 ;
        RECT 1.3350 0.6825 1.3950 0.7425 ;
        RECT 1.2300 0.4950 1.2900 0.5550 ;
        RECT 1.1250 0.1725 1.1850 0.2325 ;
        RECT 1.1250 0.8475 1.1850 0.9075 ;
        RECT 1.0200 0.4950 1.0800 0.5550 ;
        RECT 0.9150 0.3225 0.9750 0.3825 ;
        RECT 0.9150 0.7575 0.9750 0.8175 ;
        RECT 0.8100 0.4950 0.8700 0.5550 ;
        RECT 0.7050 0.1725 0.7650 0.2325 ;
        RECT 0.7050 0.6825 0.7650 0.7425 ;
        RECT 0.6000 0.4950 0.6600 0.5550 ;
        RECT 0.4950 0.3225 0.5550 0.3825 ;
        RECT 0.4950 0.8325 0.5550 0.8925 ;
        RECT 0.3900 0.4950 0.4500 0.5550 ;
        RECT 0.2850 0.1725 0.3450 0.2325 ;
        RECT 0.2850 0.6825 0.3450 0.7425 ;
        RECT 0.1800 0.4950 0.2400 0.5550 ;
        RECT 0.0750 0.2550 0.1350 0.3150 ;
        RECT 0.0750 0.7800 0.1350 0.8400 ;
        LAYER M1 ;
        RECT 3.6375 0.7125 3.7125 0.8475 ;
        RECT 3.2925 0.7125 3.6375 0.7875 ;
        RECT 3.4275 0.2100 3.5025 0.3900 ;
        RECT 3.0825 0.3150 3.4275 0.3900 ;
        RECT 3.2175 0.6600 3.2925 0.7875 ;
        RECT 2.8725 0.6600 3.2175 0.7350 ;
        RECT 3.0075 0.2100 3.0825 0.3900 ;
        RECT 2.6625 0.3150 3.0075 0.3900 ;
        RECT 2.7975 0.6600 2.8725 0.8475 ;
        RECT 2.0325 0.6600 2.7975 0.7350 ;
        RECT 2.0400 0.4725 2.7900 0.5775 ;
        RECT 2.1450 0.8100 2.6850 0.8850 ;
        RECT 2.5875 0.2100 2.6625 0.3900 ;
        RECT 2.2425 0.3150 2.5875 0.3900 ;
        RECT 2.1675 0.2100 2.2425 0.3900 ;
        RECT 1.9575 0.6600 2.0325 0.8475 ;
        RECT 1.7475 0.2100 1.8225 0.3900 ;
        RECT 1.7475 0.6750 1.8225 0.8475 ;
        RECT 0.1425 0.3150 1.7475 0.3900 ;
        RECT 0.9825 0.6750 1.7475 0.7500 ;
        RECT 0.9900 0.4725 1.7400 0.5775 ;
        RECT 0.2550 0.1650 1.6350 0.2400 ;
        RECT 0.9075 0.6750 0.9825 0.9000 ;
        RECT 0.1500 0.4725 0.9150 0.5775 ;
        RECT 0.1425 0.8250 0.9075 0.9000 ;
        RECT 0.2550 0.6750 0.7950 0.7500 ;
        RECT 0.0675 0.2250 0.1425 0.3900 ;
        RECT 0.0675 0.7500 0.1425 0.9000 ;
        LAYER VIA1 ;
        RECT 2.1900 0.8100 2.2650 0.8850 ;
        RECT 2.1675 0.2550 2.2425 0.3300 ;
        RECT 1.7475 0.2625 1.8225 0.3375 ;
        RECT 1.4325 0.1650 1.5075 0.2400 ;
        LAYER M2 ;
        RECT 2.0325 0.8100 2.3100 0.8850 ;
        RECT 2.1675 0.1125 2.2425 0.3750 ;
        RECT 1.5225 0.1125 2.1675 0.1875 ;
        RECT 1.9575 0.2625 2.0325 0.8850 ;
        RECT 1.6725 0.2625 1.9575 0.3375 ;
        RECT 1.4175 0.1125 1.5225 0.2775 ;
    END
END OAI22_0111


MACRO OAI22_1000
    CLASS CORE ;
    FOREIGN OAI22_1000 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.0500 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 0.4650 0.1125 0.8700 0.1875 ;
        RECT 0.3600 0.1125 0.4650 0.4575 ;
        VIA 0.4125 0.3825 VIA12_square ;
        END
    END ZN
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.9075 0.4125 1.0125 0.6825 ;
        RECT 0.7800 0.4125 0.9075 0.5775 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.4800 0.7125 0.9450 0.7875 ;
        VIA 0.6675 0.7500 VIA12_square ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.0675 0.5625 0.5400 0.6375 ;
        VIA 0.2625 0.6000 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.3600 0.8625 0.8250 0.9375 ;
        RECT 0.2550 0.7725 0.3600 0.9375 ;
        VIA 0.3075 0.8550 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.7950 -0.0750 1.0500 0.0750 ;
        RECT 0.6750 -0.0750 0.7950 0.1875 ;
        RECT 0.0000 -0.0750 0.6750 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.0050 0.9750 1.0500 1.1250 ;
        RECT 0.8850 0.8025 1.0050 1.1250 ;
        RECT 0.1200 0.9750 0.8850 1.1250 ;
        RECT 0.1200 0.6525 0.1500 0.7800 ;
        RECT 0.0450 0.6525 0.1200 1.1250 ;
        RECT 0.0000 0.9750 0.0450 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 0.9150 0.1575 0.9750 0.2175 ;
        RECT 0.9150 0.8325 0.9750 0.8925 ;
        RECT 0.8175 0.4875 0.8775 0.5475 ;
        RECT 0.7050 0.1200 0.7650 0.1800 ;
        RECT 0.6000 0.4575 0.6600 0.5175 ;
        RECT 0.4950 0.1575 0.5550 0.2175 ;
        RECT 0.4950 0.6300 0.5550 0.6900 ;
        RECT 0.3900 0.8400 0.4500 0.9000 ;
        RECT 0.2850 0.3000 0.3450 0.3600 ;
        RECT 0.1800 0.4950 0.2400 0.5550 ;
        RECT 0.0750 0.1650 0.1350 0.2250 ;
        RECT 0.0750 0.6825 0.1350 0.7425 ;
        LAYER M1 ;
        RECT 0.8850 0.1500 1.0050 0.3375 ;
        RECT 0.6000 0.2625 0.8850 0.3375 ;
        RECT 0.6300 0.4125 0.7050 0.8700 ;
        RECT 0.5625 0.4125 0.6300 0.5175 ;
        RECT 0.5250 0.1500 0.6000 0.3375 ;
        RECT 0.4500 0.6000 0.5550 0.7200 ;
        RECT 0.2250 0.7950 0.5550 0.9000 ;
        RECT 0.1425 0.1500 0.5250 0.2250 ;
        RECT 0.3750 0.3000 0.4500 0.7200 ;
        RECT 0.2550 0.3000 0.3750 0.4050 ;
        RECT 0.2250 0.4800 0.3000 0.6900 ;
        RECT 0.1650 0.4800 0.2250 0.5775 ;
        RECT 0.0600 0.4050 0.1650 0.5775 ;
        RECT 0.0375 0.1500 0.1425 0.2550 ;
    END
END OAI22_1000


MACRO OAI22_1010
    CLASS CORE ;
    FOREIGN OAI22_1010 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.0500 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.4500 0.6150 0.5925 0.7200 ;
        RECT 0.3750 0.3000 0.4500 0.7200 ;
        RECT 0.2625 0.3000 0.3750 0.4050 ;
        END
    END ZN
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.9075 0.4125 1.0125 0.6825 ;
        RECT 0.8175 0.4125 0.9075 0.5775 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.6675 0.4125 0.7425 0.8700 ;
        RECT 0.5625 0.4125 0.6675 0.5400 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.2250 0.4800 0.3000 0.6900 ;
        RECT 0.1650 0.4800 0.2250 0.5775 ;
        RECT 0.0600 0.3675 0.1650 0.5775 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.3600 0.8625 0.5550 0.9375 ;
        RECT 0.2550 0.7725 0.3600 0.9375 ;
        RECT 0.0900 0.8625 0.2550 0.9375 ;
        VIA 0.3075 0.8550 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.7950 -0.0750 1.0500 0.0750 ;
        RECT 0.6750 -0.0750 0.7950 0.1875 ;
        RECT 0.0000 -0.0750 0.6750 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.0050 0.9750 1.0500 1.1250 ;
        RECT 0.8850 0.7875 1.0050 1.1250 ;
        RECT 0.1200 0.9750 0.8850 1.1250 ;
        RECT 0.1200 0.6525 0.1500 0.7800 ;
        RECT 0.0450 0.6525 0.1200 1.1250 ;
        RECT 0.0000 0.9750 0.0450 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 0.9150 0.2175 0.9750 0.2775 ;
        RECT 0.9150 0.7875 0.9750 0.8475 ;
        RECT 0.8175 0.4875 0.8775 0.5475 ;
        RECT 0.7050 0.1200 0.7650 0.1800 ;
        RECT 0.6000 0.4800 0.6600 0.5400 ;
        RECT 0.4950 0.1575 0.5550 0.2175 ;
        RECT 0.4950 0.6600 0.5550 0.7200 ;
        RECT 0.3900 0.8400 0.4500 0.9000 ;
        RECT 0.2850 0.3225 0.3450 0.3825 ;
        RECT 0.1800 0.4950 0.2400 0.5550 ;
        RECT 0.0750 0.1650 0.1350 0.2250 ;
        RECT 0.0750 0.6825 0.1350 0.7425 ;
        LAYER M1 ;
        RECT 0.8925 0.1800 0.9825 0.3375 ;
        RECT 0.6000 0.2625 0.8925 0.3375 ;
        RECT 0.5250 0.1500 0.6000 0.3375 ;
        RECT 0.2250 0.7950 0.5550 0.9000 ;
        RECT 0.1425 0.1500 0.5250 0.2250 ;
        RECT 0.0375 0.1500 0.1425 0.2550 ;
    END
END OAI22_1010


MACRO OAI31_0011
    CLASS CORE ;
    FOREIGN OAI31_0011 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.8900 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 0.9825 0.7125 1.4475 0.7875 ;
        RECT 0.9825 0.2700 1.0125 0.4200 ;
        RECT 0.9075 0.2700 0.9825 0.7875 ;
        VIA 1.2525 0.7500 VIA12_square ;
        VIA 0.9600 0.3450 VIA12_square ;
        END
    END ZN
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.7475 0.4125 1.8225 0.6825 ;
        RECT 1.6575 0.4125 1.7475 0.5850 ;
        RECT 1.4475 0.4650 1.6575 0.5850 ;
        END
    END B
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.8325 0.8625 1.2975 0.9375 ;
        RECT 0.7575 0.3975 0.8325 0.9375 ;
        VIA 0.7950 0.5250 VIA12_square ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.6075 0.5475 0.6825 0.9375 ;
        RECT 0.1425 0.8625 0.6075 0.9375 ;
        VIA 0.6450 0.6900 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.1925 0.4875 1.3875 0.5625 ;
        RECT 1.1175 0.1125 1.1925 0.5625 ;
        RECT 0.4275 0.1125 1.1175 0.1875 ;
        RECT 0.3525 0.1125 0.4275 0.6375 ;
        RECT 0.0600 0.5625 0.3525 0.6375 ;
        VIA 1.2750 0.5250 VIA12_square ;
        VIA 0.1725 0.6000 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.6350 -0.0750 1.8900 0.0750 ;
        RECT 1.5150 -0.0750 1.6350 0.1875 ;
        RECT 0.0000 -0.0750 1.5150 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.8225 0.9750 1.8900 1.1250 ;
        RECT 1.7475 0.7875 1.8225 1.1250 ;
        RECT 1.4250 0.9750 1.7475 1.1250 ;
        RECT 1.3050 0.8625 1.4250 1.1250 ;
        RECT 0.1575 0.9750 1.3050 1.1250 ;
        RECT 0.0525 0.7500 0.1575 1.1250 ;
        RECT 0.0000 0.9750 0.0525 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.7550 0.2475 1.8150 0.3075 ;
        RECT 1.7550 0.8175 1.8150 0.8775 ;
        RECT 1.6500 0.4950 1.7100 0.5550 ;
        RECT 1.5450 0.1200 1.6050 0.1800 ;
        RECT 1.5450 0.7575 1.6050 0.8175 ;
        RECT 1.4475 0.4950 1.5075 0.5550 ;
        RECT 1.3350 0.2325 1.3950 0.2925 ;
        RECT 1.3350 0.8700 1.3950 0.9300 ;
        RECT 1.2300 0.4950 1.2900 0.5550 ;
        RECT 1.1250 0.3150 1.1850 0.3750 ;
        RECT 1.0200 0.4950 1.0800 0.5550 ;
        RECT 0.9150 0.1575 0.9750 0.2175 ;
        RECT 0.8100 0.4950 0.8700 0.5550 ;
        RECT 0.7050 0.3150 0.7650 0.3750 ;
        RECT 0.7050 0.8250 0.7650 0.8850 ;
        RECT 0.6000 0.4950 0.6600 0.5550 ;
        RECT 0.4950 0.1575 0.5550 0.2175 ;
        RECT 0.3900 0.4950 0.4500 0.5550 ;
        RECT 0.2850 0.3150 0.3450 0.3750 ;
        RECT 0.1725 0.4950 0.2325 0.5550 ;
        RECT 0.0750 0.1725 0.1350 0.2325 ;
        RECT 0.0750 0.7725 0.1350 0.8325 ;
        LAYER M1 ;
        RECT 1.7325 0.2250 1.8375 0.3375 ;
        RECT 1.4025 0.2625 1.7325 0.3375 ;
        RECT 1.5375 0.7125 1.6125 0.8475 ;
        RECT 1.2075 0.7125 1.5375 0.7875 ;
        RECT 1.3275 0.1500 1.4025 0.3375 ;
        RECT 1.1775 0.4725 1.3725 0.6375 ;
        RECT 0.1650 0.1500 1.3275 0.2250 ;
        RECT 0.2550 0.3000 1.2150 0.3975 ;
        RECT 1.1325 0.7125 1.2075 0.9000 ;
        RECT 0.6750 0.8025 1.1325 0.9000 ;
        RECT 1.0575 0.4725 1.1025 0.5775 ;
        RECT 0.9825 0.4725 1.0575 0.7275 ;
        RECT 0.4800 0.6525 0.9825 0.7275 ;
        RECT 0.5775 0.4725 0.8925 0.5775 ;
        RECT 0.3600 0.4950 0.4800 0.7275 ;
        RECT 0.0825 0.4725 0.2625 0.6750 ;
        RECT 0.0450 0.1500 0.1650 0.2550 ;
    END
END OAI31_0011


MACRO OAI31_0111
    CLASS CORE ;
    FOREIGN OAI31_0111 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.7800 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 0.3675 0.2700 0.6825 0.7875 ;
        VIA 0.5250 0.3525 VIA12_slot ;
        VIA 0.5250 0.7050 VIA12_slot ;
        END
    END ZN
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 3.6375 0.4125 3.7125 0.6825 ;
        RECT 3.5475 0.4125 3.6375 0.5850 ;
        RECT 2.9025 0.4650 3.5475 0.5850 ;
        END
    END B
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1425 0.4800 0.9000 0.5850 ;
        RECT 0.0675 0.3675 0.1425 0.6825 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.4025 0.5625 1.7175 0.6375 ;
        RECT 1.3275 0.4125 1.4025 0.6375 ;
        RECT 1.0125 0.4125 1.3275 0.4875 ;
        VIA 1.3650 0.5325 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 2.2425 0.5625 2.5575 0.6375 ;
        RECT 2.1675 0.4125 2.2425 0.6375 ;
        RECT 1.8525 0.4125 2.1675 0.4875 ;
        VIA 2.2050 0.5250 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 3.5250 -0.0750 3.7800 0.0750 ;
        RECT 3.4050 -0.0750 3.5250 0.1875 ;
        RECT 3.0975 -0.0750 3.4050 0.0750 ;
        RECT 2.9925 -0.0750 3.0975 0.2400 ;
        RECT 0.0000 -0.0750 2.9925 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 3.7125 0.9750 3.7800 1.1250 ;
        RECT 3.6375 0.7875 3.7125 1.1250 ;
        RECT 3.3150 0.9750 3.6375 1.1250 ;
        RECT 3.1950 0.8400 3.3150 1.1250 ;
        RECT 2.8725 0.9750 3.1950 1.1250 ;
        RECT 2.7975 0.7425 2.8725 1.1250 ;
        RECT 2.4675 0.9750 2.7975 1.1250 ;
        RECT 2.3625 0.8100 2.4675 1.1250 ;
        RECT 2.0550 0.9750 2.3625 1.1250 ;
        RECT 1.9500 0.8025 2.0550 1.1250 ;
        RECT 0.0000 0.9750 1.9500 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 3.6450 0.2400 3.7050 0.3000 ;
        RECT 3.6450 0.8175 3.7050 0.8775 ;
        RECT 3.5400 0.4950 3.6000 0.5550 ;
        RECT 3.4350 0.1200 3.4950 0.1800 ;
        RECT 3.4350 0.6825 3.4950 0.7425 ;
        RECT 3.3300 0.4950 3.3900 0.5550 ;
        RECT 3.2250 0.2925 3.2850 0.3525 ;
        RECT 3.2250 0.8475 3.2850 0.9075 ;
        RECT 3.1200 0.4950 3.1800 0.5550 ;
        RECT 3.0150 0.1575 3.0750 0.2175 ;
        RECT 3.0150 0.6825 3.0750 0.7425 ;
        RECT 2.9100 0.4950 2.9700 0.5550 ;
        RECT 2.8050 0.2475 2.8650 0.3075 ;
        RECT 2.8050 0.7725 2.8650 0.8325 ;
        RECT 2.7000 0.4950 2.7600 0.5550 ;
        RECT 2.5950 0.3225 2.6550 0.3825 ;
        RECT 2.5950 0.6675 2.6550 0.7275 ;
        RECT 2.4900 0.4950 2.5500 0.5550 ;
        RECT 2.3850 0.1575 2.4450 0.2175 ;
        RECT 2.3850 0.8325 2.4450 0.8925 ;
        RECT 2.2800 0.4950 2.3400 0.5550 ;
        RECT 2.1750 0.3225 2.2350 0.3825 ;
        RECT 2.1750 0.6675 2.2350 0.7275 ;
        RECT 2.0700 0.4950 2.1300 0.5550 ;
        RECT 1.9650 0.1575 2.0250 0.2175 ;
        RECT 1.9650 0.8325 2.0250 0.8925 ;
        RECT 1.7550 0.1575 1.8150 0.2175 ;
        RECT 1.7550 0.8325 1.8150 0.8925 ;
        RECT 1.6500 0.4950 1.7100 0.5550 ;
        RECT 1.5450 0.3225 1.6050 0.3825 ;
        RECT 1.5450 0.6675 1.6050 0.7275 ;
        RECT 1.4400 0.4950 1.5000 0.5550 ;
        RECT 1.3350 0.1575 1.3950 0.2175 ;
        RECT 1.3350 0.8325 1.3950 0.8925 ;
        RECT 1.2300 0.4950 1.2900 0.5550 ;
        RECT 1.1250 0.3225 1.1850 0.3825 ;
        RECT 1.1250 0.6675 1.1850 0.7275 ;
        RECT 1.0200 0.4950 1.0800 0.5550 ;
        RECT 0.9150 0.1575 0.9750 0.2175 ;
        RECT 0.9150 0.8325 0.9750 0.8925 ;
        RECT 0.8100 0.4950 0.8700 0.5550 ;
        RECT 0.7050 0.3225 0.7650 0.3825 ;
        RECT 0.7050 0.6750 0.7650 0.7350 ;
        RECT 0.6000 0.4950 0.6600 0.5550 ;
        RECT 0.4950 0.1575 0.5550 0.2175 ;
        RECT 0.4950 0.8325 0.5550 0.8925 ;
        RECT 0.3900 0.4950 0.4500 0.5550 ;
        RECT 0.2850 0.3225 0.3450 0.3825 ;
        RECT 0.2850 0.6750 0.3450 0.7350 ;
        RECT 0.1800 0.4950 0.2400 0.5550 ;
        RECT 0.0750 0.1800 0.1350 0.2400 ;
        RECT 0.0750 0.8100 0.1350 0.8700 ;
        LAYER M1 ;
        RECT 3.6225 0.2175 3.7275 0.3375 ;
        RECT 3.3225 0.2625 3.6225 0.3375 ;
        RECT 2.9625 0.6600 3.5175 0.7650 ;
        RECT 3.1875 0.2625 3.3225 0.3900 ;
        RECT 2.8725 0.3150 3.1875 0.3900 ;
        RECT 2.7975 0.1500 2.8725 0.3900 ;
        RECT 0.1575 0.1500 2.7975 0.2250 ;
        RECT 2.0400 0.4800 2.7900 0.5775 ;
        RECT 0.2550 0.3000 2.7225 0.4050 ;
        RECT 1.8900 0.6525 2.6850 0.7275 ;
        RECT 1.8150 0.6525 1.8900 0.7350 ;
        RECT 0.1575 0.8250 1.8450 0.9000 ;
        RECT 1.0950 0.6600 1.8150 0.7350 ;
        RECT 0.9900 0.4800 1.7400 0.5850 ;
        RECT 0.2550 0.6600 0.7950 0.7500 ;
        RECT 0.0525 0.1500 0.1575 0.2625 ;
        RECT 0.0525 0.7875 0.1575 0.9000 ;
        LAYER VIA1 ;
        RECT 3.0075 0.6750 3.0825 0.7500 ;
        RECT 2.6025 0.3150 2.6775 0.3900 ;
        LAYER M2 ;
        RECT 2.7975 0.6750 3.1575 0.7500 ;
        RECT 2.7225 0.3150 2.7975 0.7500 ;
        RECT 2.5275 0.3150 2.7225 0.3900 ;
    END
END OAI31_0111


MACRO OAI31_1000
    CLASS CORE ;
    FOREIGN OAI31_1000 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.2600 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.9450 0.6675 0.9975 0.9000 ;
        RECT 0.8700 0.3075 0.9450 0.9000 ;
        RECT 0.2550 0.3075 0.8700 0.3825 ;
        RECT 0.6825 0.7800 0.8700 0.9000 ;
        END
    END ZN
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.1175 0.3675 1.1925 0.6825 ;
        RECT 1.0200 0.4500 1.1175 0.5700 ;
        END
    END B
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.5925 0.4575 0.7725 0.7050 ;
        RECT 0.4875 0.6225 0.5925 0.8325 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.3900 0.4725 0.4800 0.5475 ;
        RECT 0.3150 0.4725 0.3900 0.8325 ;
        RECT 0.2775 0.6675 0.3150 0.8325 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1425 0.4575 0.2400 0.5775 ;
        RECT 0.0675 0.3675 0.1425 0.6825 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.2150 -0.0750 1.2600 0.0750 ;
        RECT 1.1100 -0.0750 1.2150 0.2475 ;
        RECT 0.0000 -0.0750 1.1100 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.2075 0.9750 1.2600 1.1250 ;
        RECT 1.1025 0.7875 1.2075 1.1250 ;
        RECT 0.1650 0.9750 1.1025 1.1250 ;
        RECT 0.0450 0.8175 0.1650 1.1250 ;
        RECT 0.0000 0.9750 0.0450 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.1250 0.1575 1.1850 0.2175 ;
        RECT 1.1250 0.8175 1.1850 0.8775 ;
        RECT 1.0200 0.4800 1.0800 0.5400 ;
        RECT 0.9150 0.1575 0.9750 0.2175 ;
        RECT 0.9150 0.8175 0.9750 0.8775 ;
        RECT 0.7050 0.3075 0.7650 0.3675 ;
        RECT 0.7050 0.8175 0.7650 0.8775 ;
        RECT 0.6000 0.4875 0.6600 0.5475 ;
        RECT 0.4950 0.1575 0.5550 0.2175 ;
        RECT 0.3900 0.4800 0.4500 0.5400 ;
        RECT 0.2850 0.3075 0.3450 0.3675 ;
        RECT 0.1800 0.4875 0.2400 0.5475 ;
        RECT 0.0750 0.1725 0.1350 0.2325 ;
        RECT 0.0750 0.8325 0.1350 0.8925 ;
        LAYER M1 ;
        RECT 0.1575 0.1500 1.0050 0.2250 ;
        RECT 0.0525 0.1500 0.1575 0.2550 ;
    END
END OAI31_1000


MACRO OAI31_1010
    CLASS CORE ;
    FOREIGN OAI31_1010 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.2600 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.9450 0.6675 0.9825 0.9000 ;
        RECT 0.8700 0.3075 0.9450 0.9000 ;
        RECT 0.2550 0.3075 0.8700 0.3825 ;
        RECT 0.7050 0.7800 0.8700 0.9000 ;
        END
    END ZN
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.1175 0.3675 1.1925 0.6825 ;
        RECT 1.0200 0.4500 1.1175 0.5700 ;
        END
    END B
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.5925 0.4575 0.7725 0.7050 ;
        RECT 0.4875 0.6225 0.5925 0.8325 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.3900 0.4725 0.4800 0.5475 ;
        RECT 0.3150 0.4725 0.3900 0.8325 ;
        RECT 0.2775 0.6675 0.3150 0.8325 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1425 0.4575 0.2400 0.5775 ;
        RECT 0.0675 0.3675 0.1425 0.6825 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.2150 -0.0750 1.2600 0.0750 ;
        RECT 1.1100 -0.0750 1.2150 0.2475 ;
        RECT 0.0000 -0.0750 1.1100 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.2075 0.9750 1.2600 1.1250 ;
        RECT 1.1025 0.7875 1.2075 1.1250 ;
        RECT 0.1650 0.9750 1.1025 1.1250 ;
        RECT 0.0450 0.8175 0.1650 1.1250 ;
        RECT 0.0000 0.9750 0.0450 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.1250 0.1575 1.1850 0.2175 ;
        RECT 1.1250 0.8175 1.1850 0.8775 ;
        RECT 1.0200 0.4800 1.0800 0.5400 ;
        RECT 0.9150 0.1575 0.9750 0.2175 ;
        RECT 0.9150 0.8100 0.9750 0.8700 ;
        RECT 0.7050 0.3075 0.7650 0.3675 ;
        RECT 0.7050 0.8100 0.7650 0.8700 ;
        RECT 0.6000 0.4875 0.6600 0.5475 ;
        RECT 0.4950 0.1575 0.5550 0.2175 ;
        RECT 0.3900 0.4800 0.4500 0.5400 ;
        RECT 0.2850 0.3075 0.3450 0.3675 ;
        RECT 0.1800 0.4875 0.2400 0.5475 ;
        RECT 0.0750 0.1725 0.1350 0.2325 ;
        RECT 0.0750 0.8325 0.1350 0.8925 ;
        LAYER M1 ;
        RECT 0.1575 0.1500 1.0050 0.2250 ;
        RECT 0.0525 0.1500 0.1575 0.2550 ;
    END
END OAI31_1010


MACRO OAI32_0011
    CLASS CORE ;
    FOREIGN OAI32_0011 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.3100 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 1.5300 0.7950 1.6800 0.9375 ;
        RECT 1.2150 0.8625 1.5300 0.9375 ;
        RECT 1.1400 0.2625 1.2150 0.9375 ;
        RECT 0.8250 0.2625 1.1400 0.3375 ;
        VIA 1.6050 0.8475 VIA12_square ;
        VIA 1.1775 0.8475 VIA12_square ;
        VIA 1.1775 0.3450 VIA12_square ;
        END
    END ZN
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.8750 0.8625 2.1900 0.9375 ;
        RECT 1.8000 0.4125 1.8750 0.9375 ;
        RECT 1.4850 0.4125 1.8000 0.4875 ;
        VIA 1.8375 0.5250 VIA12_square ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 2.0700 0.4125 2.2425 0.7350 ;
        RECT 1.5525 0.6600 2.0700 0.7350 ;
        RECT 1.4775 0.4575 1.5525 0.7350 ;
        RECT 1.4400 0.4575 1.4775 0.5775 ;
        END
    END B1
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.8100 0.4125 1.0125 0.4875 ;
        RECT 0.6600 0.4125 0.8100 0.5775 ;
        RECT 0.5475 0.4125 0.6600 0.4875 ;
        VIA 0.7350 0.5250 VIA12_square ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.9075 0.6150 1.0125 0.7875 ;
        RECT 0.4425 0.7125 0.9075 0.7875 ;
        VIA 0.9600 0.6975 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.2900 0.1125 1.3650 0.6375 ;
        RECT 0.4275 0.1125 1.2900 0.1875 ;
        RECT 0.3525 0.1125 0.4275 0.6375 ;
        RECT 0.0975 0.5625 0.3525 0.6375 ;
        VIA 1.3275 0.5550 VIA12_square ;
        VIA 0.2100 0.6000 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 2.0550 -0.0750 2.3100 0.0750 ;
        RECT 1.9350 -0.0750 2.0550 0.1875 ;
        RECT 1.6275 -0.0750 1.9350 0.0750 ;
        RECT 1.5225 -0.0750 1.6275 0.2325 ;
        RECT 0.0000 -0.0750 1.5225 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 2.2650 0.9750 2.3100 1.1250 ;
        RECT 2.1450 0.8100 2.2650 1.1250 ;
        RECT 1.4025 0.9750 2.1450 1.1250 ;
        RECT 1.3275 0.7725 1.4025 1.1250 ;
        RECT 0.1575 0.9750 1.3275 1.1250 ;
        RECT 0.0525 0.7500 0.1575 1.1250 ;
        RECT 0.0000 0.9750 0.0525 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 2.1750 0.2250 2.2350 0.2850 ;
        RECT 2.1750 0.8175 2.2350 0.8775 ;
        RECT 2.0700 0.4950 2.1300 0.5550 ;
        RECT 1.9650 0.1200 2.0250 0.1800 ;
        RECT 1.8600 0.4950 1.9200 0.5550 ;
        RECT 1.7550 0.2925 1.8150 0.3525 ;
        RECT 1.7550 0.8250 1.8150 0.8850 ;
        RECT 1.6500 0.4950 1.7100 0.5550 ;
        RECT 1.5450 0.1500 1.6050 0.2100 ;
        RECT 1.4400 0.4875 1.5000 0.5475 ;
        RECT 1.3350 0.1575 1.3950 0.2175 ;
        RECT 1.3350 0.8025 1.3950 0.8625 ;
        RECT 1.2300 0.4875 1.2900 0.5475 ;
        RECT 1.1250 0.3150 1.1850 0.3750 ;
        RECT 1.0200 0.4950 1.0800 0.5550 ;
        RECT 0.9150 0.1575 0.9750 0.2175 ;
        RECT 0.8100 0.4950 0.8700 0.5550 ;
        RECT 0.7050 0.3225 0.7650 0.3825 ;
        RECT 0.7050 0.8250 0.7650 0.8850 ;
        RECT 0.6000 0.4950 0.6600 0.5550 ;
        RECT 0.4950 0.1575 0.5550 0.2175 ;
        RECT 0.3900 0.4950 0.4500 0.5550 ;
        RECT 0.2850 0.3225 0.3450 0.3825 ;
        RECT 0.1800 0.4950 0.2400 0.5550 ;
        RECT 0.0750 0.2250 0.1350 0.2850 ;
        RECT 0.0750 0.7725 0.1350 0.8325 ;
        LAYER M1 ;
        RECT 2.1525 0.1950 2.2575 0.3375 ;
        RECT 1.8525 0.2625 2.1525 0.3375 ;
        RECT 1.5075 0.8100 2.0025 0.9000 ;
        RECT 1.6275 0.4725 1.9425 0.5775 ;
        RECT 1.7175 0.2625 1.8525 0.3825 ;
        RECT 1.4400 0.3075 1.7175 0.3825 ;
        RECT 1.3650 0.1500 1.4400 0.3825 ;
        RECT 0.1500 0.1500 1.3650 0.2250 ;
        RECT 1.1775 0.4725 1.3650 0.6675 ;
        RECT 0.2550 0.3000 1.2600 0.3975 ;
        RECT 1.1025 0.7950 1.2525 0.9000 ;
        RECT 1.0425 0.4725 1.1025 0.5775 ;
        RECT 0.6750 0.8100 1.1025 0.9000 ;
        RECT 0.9675 0.4725 1.0425 0.7350 ;
        RECT 0.5025 0.6600 0.9675 0.7350 ;
        RECT 0.5775 0.4725 0.8925 0.5775 ;
        RECT 0.4275 0.4725 0.5025 0.7350 ;
        RECT 0.3675 0.4725 0.4275 0.5775 ;
        RECT 0.0975 0.4725 0.2925 0.6750 ;
        RECT 0.0600 0.1500 0.1500 0.3150 ;
    END
END OAI32_0011


MACRO OAI32_0111
    CLASS CORE ;
    FOREIGN OAI32_0111 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.5200 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 1.8375 0.2625 2.1525 0.7500 ;
        VIA 1.9950 0.3450 VIA12_slot ;
        VIA 1.9950 0.6675 VIA12_slot ;
        END
    END ZN
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.8775 0.7125 1.3425 0.7875 ;
        VIA 0.9900 0.7500 VIA12_square ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.9750 0.5625 1.4400 0.6375 ;
        VIA 1.1550 0.6000 VIA12_square ;
        END
    END B1
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.7275 0.2625 1.1775 0.3375 ;
        RECT 0.7275 0.5025 0.7575 0.6075 ;
        RECT 0.6525 0.2625 0.7275 0.6075 ;
        VIA 0.6900 0.5250 VIA12_square ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.0675 0.7125 0.5325 0.7875 ;
        VIA 0.4200 0.7500 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.5025 0.5325 0.5775 0.6375 ;
        RECT 0.1125 0.5625 0.5025 0.6375 ;
        VIA 0.2400 0.6000 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 2.4525 -0.0750 2.5200 0.0750 ;
        RECT 2.3775 -0.0750 2.4525 0.3150 ;
        RECT 2.0550 -0.0750 2.3775 0.0750 ;
        RECT 1.9350 -0.0750 2.0550 0.1950 ;
        RECT 1.6350 -0.0750 1.9350 0.0750 ;
        RECT 1.5150 -0.0750 1.6350 0.1875 ;
        RECT 1.0050 -0.0750 1.5150 0.0750 ;
        RECT 0.8850 -0.0750 1.0050 0.1875 ;
        RECT 0.0000 -0.0750 0.8850 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 2.4525 0.9750 2.5200 1.1250 ;
        RECT 2.3775 0.6375 2.4525 1.1250 ;
        RECT 2.0325 0.9750 2.3775 1.1250 ;
        RECT 1.9575 0.8175 2.0325 1.1250 ;
        RECT 1.6350 0.9750 1.9575 1.1250 ;
        RECT 1.5150 0.8175 1.6350 1.1250 ;
        RECT 1.2075 0.9750 1.5150 1.1250 ;
        RECT 1.1025 0.7950 1.2075 1.1250 ;
        RECT 0.1425 0.9750 1.1025 1.1250 ;
        RECT 0.0675 0.7950 0.1425 1.1250 ;
        RECT 0.0000 0.9750 0.0675 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 2.3850 0.2250 2.4450 0.2850 ;
        RECT 2.3850 0.6675 2.4450 0.7275 ;
        RECT 2.3850 0.8325 2.4450 0.8925 ;
        RECT 2.2800 0.4650 2.3400 0.5250 ;
        RECT 2.1750 0.2250 2.2350 0.2850 ;
        RECT 2.1750 0.7200 2.2350 0.7800 ;
        RECT 2.0700 0.4650 2.1300 0.5250 ;
        RECT 1.9650 0.1275 2.0250 0.1875 ;
        RECT 1.9650 0.8475 2.0250 0.9075 ;
        RECT 1.8600 0.4650 1.9200 0.5250 ;
        RECT 1.7550 0.2250 1.8150 0.2850 ;
        RECT 1.7550 0.7200 1.8150 0.7800 ;
        RECT 1.6500 0.4650 1.7100 0.5250 ;
        RECT 1.5450 0.1275 1.6050 0.1875 ;
        RECT 1.5450 0.8250 1.6050 0.8850 ;
        RECT 1.4400 0.4650 1.5000 0.5250 ;
        RECT 1.3350 0.2250 1.3950 0.2850 ;
        RECT 1.3350 0.7575 1.3950 0.8175 ;
        RECT 1.1250 0.1575 1.1850 0.2175 ;
        RECT 1.1250 0.8250 1.1850 0.8850 ;
        RECT 1.0200 0.4650 1.0800 0.5250 ;
        RECT 0.9150 0.1275 0.9750 0.1875 ;
        RECT 0.8175 0.4950 0.8775 0.5550 ;
        RECT 0.7050 0.1575 0.7650 0.2175 ;
        RECT 0.7050 0.8175 0.7650 0.8775 ;
        RECT 0.6000 0.4950 0.6600 0.5550 ;
        RECT 0.4950 0.3075 0.5550 0.3675 ;
        RECT 0.3900 0.4950 0.4500 0.5550 ;
        RECT 0.2850 0.1575 0.3450 0.2175 ;
        RECT 0.1800 0.4950 0.2400 0.5550 ;
        RECT 0.0750 0.1800 0.1350 0.2400 ;
        RECT 0.0750 0.8325 0.1350 0.8925 ;
        LAYER M1 ;
        RECT 1.6575 0.4575 2.3700 0.5325 ;
        RECT 2.1525 0.1950 2.2575 0.3825 ;
        RECT 2.1675 0.6225 2.2425 0.8325 ;
        RECT 1.8225 0.6225 2.1675 0.7125 ;
        RECT 1.8375 0.2925 2.1525 0.3825 ;
        RECT 1.7325 0.1950 1.8375 0.3825 ;
        RECT 1.7475 0.6225 1.8225 0.8325 ;
        RECT 1.5825 0.2625 1.6575 0.7125 ;
        RECT 1.4175 0.2625 1.5825 0.3375 ;
        RECT 1.4025 0.6375 1.5825 0.7125 ;
        RECT 1.2825 0.4125 1.5000 0.5625 ;
        RECT 1.3125 0.1950 1.4175 0.3375 ;
        RECT 1.3275 0.6375 1.4025 0.8700 ;
        RECT 1.0950 0.1500 1.2150 0.3375 ;
        RECT 1.1025 0.4125 1.2075 0.6825 ;
        RECT 0.9750 0.4125 1.1025 0.5250 ;
        RECT 0.8100 0.2625 1.0950 0.3375 ;
        RECT 0.9525 0.6000 1.0275 0.8475 ;
        RECT 0.9000 0.6000 0.9525 0.6750 ;
        RECT 0.8175 0.4650 0.9000 0.6750 ;
        RECT 0.5625 0.7500 0.8475 0.9000 ;
        RECT 0.7350 0.1500 0.8100 0.3375 ;
        RECT 0.5475 0.4500 0.7425 0.6150 ;
        RECT 0.2550 0.1500 0.7350 0.2250 ;
        RECT 0.1500 0.3000 0.6075 0.3750 ;
        RECT 0.3675 0.4725 0.4725 0.8325 ;
        RECT 0.2175 0.4500 0.2925 0.8400 ;
        RECT 0.1800 0.4500 0.2175 0.6825 ;
        RECT 0.0450 0.1500 0.1500 0.3750 ;
        LAYER VIA1 ;
        RECT 1.3725 0.4125 1.4475 0.4875 ;
        RECT 0.6675 0.8025 0.7425 0.8775 ;
        RECT 0.4125 0.3000 0.4875 0.3750 ;
        LAYER M2 ;
        RECT 1.5600 0.4125 1.6350 0.9375 ;
        RECT 1.4025 0.4125 1.5600 0.4875 ;
        RECT 0.7575 0.8625 1.5600 0.9375 ;
        RECT 1.3275 0.1125 1.4025 0.4875 ;
        RECT 0.5475 0.1125 1.3275 0.1875 ;
        RECT 0.6525 0.7500 0.7575 0.9375 ;
        RECT 0.4725 0.1125 0.5475 0.3750 ;
        RECT 0.3525 0.3000 0.4725 0.3750 ;
    END
END OAI32_0111


MACRO OAI32_1000
    CLASS CORE ;
    FOREIGN OAI32_1000 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.4700 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 0.7725 0.7125 0.8925 0.7875 ;
        RECT 0.6975 0.1125 0.7725 0.7875 ;
        RECT 0.2325 0.1125 0.6975 0.1875 ;
        VIA 0.7800 0.7500 VIA12_square ;
        VIA 0.7350 0.3375 VIA12_square ;
        END
    END ZN
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.0725 0.7425 1.1775 0.9375 ;
        RECT 0.6075 0.8625 1.0725 0.9375 ;
        VIA 1.1250 0.8175 VIA12_square ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.3125 0.4125 1.4175 0.6825 ;
        RECT 1.1850 0.4125 1.3125 0.5475 ;
        END
    END B1
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.9225 0.1125 1.3875 0.1875 ;
        RECT 0.9225 0.4725 0.9525 0.6375 ;
        RECT 0.8475 0.1125 0.9225 0.6375 ;
        VIA 0.9000 0.5550 VIA12_square ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.1125 0.7125 0.5775 0.7875 ;
        VIA 0.4200 0.7500 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.1125 0.5625 0.5775 0.6375 ;
        VIA 0.2400 0.6000 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.2150 -0.0750 1.4700 0.0750 ;
        RECT 1.0950 -0.0750 1.2150 0.1875 ;
        RECT 0.0000 -0.0750 1.0950 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.4175 0.9750 1.4700 1.1250 ;
        RECT 1.3125 0.7950 1.4175 1.1250 ;
        RECT 0.1425 0.9750 1.3125 1.1250 ;
        RECT 0.0675 0.7950 0.1425 1.1250 ;
        RECT 0.0000 0.9750 0.0675 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.3350 0.1575 1.3950 0.2175 ;
        RECT 1.3350 0.8250 1.3950 0.8850 ;
        RECT 1.2300 0.4800 1.2900 0.5400 ;
        RECT 1.1250 0.1275 1.1850 0.1875 ;
        RECT 1.0275 0.4950 1.0875 0.5550 ;
        RECT 0.9150 0.1575 0.9750 0.2175 ;
        RECT 0.9150 0.8175 0.9750 0.8775 ;
        RECT 0.7050 0.1575 0.7650 0.2175 ;
        RECT 0.7050 0.8175 0.7650 0.8775 ;
        RECT 0.6000 0.4950 0.6600 0.5550 ;
        RECT 0.4950 0.3075 0.5550 0.3675 ;
        RECT 0.3900 0.4950 0.4500 0.5550 ;
        RECT 0.2850 0.1575 0.3450 0.2175 ;
        RECT 0.1800 0.4950 0.2400 0.5550 ;
        RECT 0.0750 0.1800 0.1350 0.2400 ;
        RECT 0.0750 0.8325 0.1350 0.8925 ;
        LAYER M1 ;
        RECT 1.3050 0.1500 1.4250 0.3375 ;
        RECT 1.0200 0.2625 1.3050 0.3375 ;
        RECT 1.1100 0.6450 1.1775 0.9000 ;
        RECT 1.0725 0.4650 1.1100 0.9000 ;
        RECT 1.0275 0.4650 1.0725 0.7200 ;
        RECT 0.9450 0.1500 1.0200 0.3375 ;
        RECT 0.8925 0.7950 0.9975 0.9000 ;
        RECT 0.8475 0.4725 0.9525 0.6375 ;
        RECT 0.2550 0.1500 0.9450 0.2250 ;
        RECT 0.6600 0.7125 0.8925 0.9000 ;
        RECT 0.5625 0.4725 0.8475 0.5925 ;
        RECT 0.1500 0.3000 0.8175 0.3750 ;
        RECT 0.3675 0.4725 0.4725 0.8325 ;
        RECT 0.2175 0.4500 0.2925 0.8400 ;
        RECT 0.1800 0.4500 0.2175 0.6825 ;
        RECT 0.0450 0.1500 0.1500 0.3750 ;
    END
END OAI32_1000


MACRO OAI32_1010
    CLASS CORE ;
    FOREIGN OAI32_1010 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.4700 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 0.7725 0.7125 0.8925 0.7875 ;
        RECT 0.6975 0.1125 0.7725 0.7875 ;
        RECT 0.2325 0.1125 0.6975 0.1875 ;
        VIA 0.7800 0.7500 VIA12_square ;
        VIA 0.7350 0.3375 VIA12_square ;
        END
    END ZN
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.0725 0.7425 1.1775 0.9375 ;
        RECT 0.6075 0.8625 1.0725 0.9375 ;
        VIA 1.1250 0.8175 VIA12_square ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.3125 0.4125 1.4175 0.6825 ;
        RECT 1.1850 0.4125 1.3125 0.5475 ;
        END
    END B1
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.9225 0.1125 1.3875 0.1875 ;
        RECT 0.9225 0.4725 0.9525 0.6375 ;
        RECT 0.8475 0.1125 0.9225 0.6375 ;
        VIA 0.9000 0.5550 VIA12_square ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.1125 0.7125 0.5775 0.7875 ;
        VIA 0.4200 0.7500 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.1125 0.5625 0.5775 0.6375 ;
        VIA 0.2400 0.6000 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.2150 -0.0750 1.4700 0.0750 ;
        RECT 1.0950 -0.0750 1.2150 0.1875 ;
        RECT 0.0000 -0.0750 1.0950 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.4175 0.9750 1.4700 1.1250 ;
        RECT 1.3125 0.7950 1.4175 1.1250 ;
        RECT 0.1425 0.9750 1.3125 1.1250 ;
        RECT 0.0675 0.7950 0.1425 1.1250 ;
        RECT 0.0000 0.9750 0.0675 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.3350 0.1575 1.3950 0.2175 ;
        RECT 1.3350 0.8250 1.3950 0.8850 ;
        RECT 1.2300 0.4800 1.2900 0.5400 ;
        RECT 1.1250 0.1275 1.1850 0.1875 ;
        RECT 1.0275 0.4950 1.0875 0.5550 ;
        RECT 0.9150 0.1575 0.9750 0.2175 ;
        RECT 0.9150 0.8175 0.9750 0.8775 ;
        RECT 0.7050 0.1575 0.7650 0.2175 ;
        RECT 0.7050 0.8175 0.7650 0.8775 ;
        RECT 0.6000 0.4950 0.6600 0.5550 ;
        RECT 0.4950 0.3075 0.5550 0.3675 ;
        RECT 0.3900 0.4950 0.4500 0.5550 ;
        RECT 0.2850 0.1575 0.3450 0.2175 ;
        RECT 0.1800 0.4950 0.2400 0.5550 ;
        RECT 0.0750 0.1800 0.1350 0.2400 ;
        RECT 0.0750 0.8325 0.1350 0.8925 ;
        LAYER M1 ;
        RECT 1.3050 0.1500 1.4250 0.3375 ;
        RECT 1.0200 0.2625 1.3050 0.3375 ;
        RECT 1.1100 0.6450 1.1775 0.9000 ;
        RECT 1.0725 0.4650 1.1100 0.9000 ;
        RECT 1.0275 0.4650 1.0725 0.7200 ;
        RECT 0.9450 0.1500 1.0200 0.3375 ;
        RECT 0.8925 0.7950 0.9975 0.9000 ;
        RECT 0.8475 0.4725 0.9525 0.6375 ;
        RECT 0.2550 0.1500 0.9450 0.2250 ;
        RECT 0.6600 0.7125 0.8925 0.9000 ;
        RECT 0.5625 0.4725 0.8475 0.5925 ;
        RECT 0.1500 0.3000 0.8175 0.3750 ;
        RECT 0.3675 0.4725 0.4725 0.8325 ;
        RECT 0.2175 0.4500 0.2925 0.8400 ;
        RECT 0.1800 0.4500 0.2175 0.6825 ;
        RECT 0.0450 0.1500 0.1500 0.3750 ;
    END
END OAI32_1010


MACRO OAI33_0011
    CLASS CORE ;
    FOREIGN OAI33_0011 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.7300 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 1.5375 0.7950 1.6875 0.9375 ;
        RECT 1.2150 0.8625 1.5375 0.9375 ;
        RECT 1.1400 0.2625 1.2150 0.9375 ;
        RECT 0.8250 0.2625 1.1400 0.3375 ;
        VIA 1.6125 0.8475 VIA12_square ;
        VIA 1.1775 0.8475 VIA12_square ;
        VIA 1.1775 0.3450 VIA12_square ;
        END
    END ZN
    PIN B3
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.9650 0.5625 2.1975 0.6375 ;
        RECT 1.8600 0.4500 1.9650 0.6375 ;
        RECT 1.7325 0.5625 1.8600 0.6375 ;
        VIA 1.9125 0.5250 VIA12_square ;
        END
    END B3
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.8525 0.7125 2.3175 0.7875 ;
        VIA 2.2050 0.7500 VIA12_square ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 2.1525 0.4125 2.6475 0.4875 ;
        RECT 2.0775 0.2625 2.1525 0.4875 ;
        RECT 1.6125 0.2625 2.0775 0.3375 ;
        RECT 1.5375 0.2625 1.6125 0.6375 ;
        RECT 1.4775 0.4875 1.5375 0.6375 ;
        VIA 2.5350 0.4500 VIA12_square ;
        VIA 1.5300 0.5625 VIA12_square ;
        END
    END B1
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.8100 0.4125 1.0125 0.4875 ;
        RECT 0.6600 0.4125 0.8100 0.5775 ;
        RECT 0.5475 0.4125 0.6600 0.4875 ;
        VIA 0.7350 0.5250 VIA12_square ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.9075 0.6150 1.0125 0.7875 ;
        RECT 0.4425 0.7125 0.9075 0.7875 ;
        VIA 0.9600 0.6975 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.2900 0.1125 1.3650 0.6375 ;
        RECT 0.4275 0.1125 1.2900 0.1875 ;
        RECT 0.3525 0.1125 0.4275 0.6375 ;
        RECT 0.0975 0.5625 0.3525 0.6375 ;
        VIA 1.3275 0.5550 VIA12_square ;
        VIA 0.2100 0.6000 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 2.4750 -0.0750 2.7300 0.0750 ;
        RECT 2.3550 -0.0750 2.4750 0.1875 ;
        RECT 2.0475 -0.0750 2.3550 0.0750 ;
        RECT 1.9425 -0.0750 2.0475 0.2325 ;
        RECT 1.6275 -0.0750 1.9425 0.0750 ;
        RECT 1.5225 -0.0750 1.6275 0.2325 ;
        RECT 0.0000 -0.0750 1.5225 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 2.6775 0.9750 2.7300 1.1250 ;
        RECT 2.5725 0.7500 2.6775 1.1250 ;
        RECT 1.4025 0.9750 2.5725 1.1250 ;
        RECT 1.3275 0.7725 1.4025 1.1250 ;
        RECT 0.1575 0.9750 1.3275 1.1250 ;
        RECT 0.0525 0.7500 0.1575 1.1250 ;
        RECT 0.0000 0.9750 0.0525 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 2.5950 0.2250 2.6550 0.2850 ;
        RECT 2.5950 0.7725 2.6550 0.8325 ;
        RECT 2.4900 0.4950 2.5500 0.5550 ;
        RECT 2.3850 0.1200 2.4450 0.1800 ;
        RECT 2.2800 0.4950 2.3400 0.5550 ;
        RECT 2.1750 0.2925 2.2350 0.3525 ;
        RECT 2.0700 0.4950 2.1300 0.5550 ;
        RECT 1.9650 0.1500 2.0250 0.2100 ;
        RECT 1.9650 0.8250 2.0250 0.8850 ;
        RECT 1.8600 0.4950 1.9200 0.5550 ;
        RECT 1.7550 0.3150 1.8150 0.3750 ;
        RECT 1.6575 0.4950 1.7175 0.5550 ;
        RECT 1.5450 0.1500 1.6050 0.2100 ;
        RECT 1.4400 0.4875 1.5000 0.5475 ;
        RECT 1.3350 0.1575 1.3950 0.2175 ;
        RECT 1.3350 0.8025 1.3950 0.8625 ;
        RECT 1.2300 0.4875 1.2900 0.5475 ;
        RECT 1.1250 0.3150 1.1850 0.3750 ;
        RECT 1.0200 0.4950 1.0800 0.5550 ;
        RECT 0.9150 0.1575 0.9750 0.2175 ;
        RECT 0.8100 0.4950 0.8700 0.5550 ;
        RECT 0.7050 0.3225 0.7650 0.3825 ;
        RECT 0.7050 0.8250 0.7650 0.8850 ;
        RECT 0.6000 0.4950 0.6600 0.5550 ;
        RECT 0.4950 0.1575 0.5550 0.2175 ;
        RECT 0.3900 0.4950 0.4500 0.5550 ;
        RECT 0.2850 0.3225 0.3450 0.3825 ;
        RECT 0.1800 0.4950 0.2400 0.5550 ;
        RECT 0.0750 0.2250 0.1350 0.2850 ;
        RECT 0.0750 0.7725 0.1350 0.8325 ;
        LAYER M1 ;
        RECT 2.5650 0.1950 2.6850 0.3375 ;
        RECT 2.4525 0.4125 2.6775 0.6300 ;
        RECT 2.2650 0.2625 2.5650 0.3375 ;
        RECT 2.3025 0.4725 2.3625 0.5775 ;
        RECT 2.2275 0.4725 2.3025 0.8325 ;
        RECT 2.1450 0.2625 2.2650 0.3825 ;
        RECT 2.1600 0.6600 2.2275 0.8325 ;
        RECT 1.7625 0.6600 2.1600 0.7350 ;
        RECT 1.8375 0.4725 2.1525 0.5775 ;
        RECT 1.4400 0.3075 2.1450 0.3825 ;
        RECT 1.5075 0.8100 2.0550 0.9000 ;
        RECT 1.6875 0.4650 1.7625 0.7350 ;
        RECT 1.6575 0.4650 1.6875 0.5850 ;
        RECT 1.4775 0.4575 1.5825 0.7200 ;
        RECT 1.4400 0.4575 1.4775 0.5925 ;
        RECT 1.3650 0.1500 1.4400 0.3825 ;
        RECT 0.1500 0.1500 1.3650 0.2250 ;
        RECT 1.1775 0.4725 1.3650 0.6675 ;
        RECT 0.2550 0.3000 1.2600 0.3975 ;
        RECT 1.1025 0.7950 1.2525 0.9000 ;
        RECT 1.0425 0.4725 1.1025 0.5775 ;
        RECT 0.6750 0.8100 1.1025 0.9000 ;
        RECT 0.9675 0.4725 1.0425 0.7350 ;
        RECT 0.5025 0.6600 0.9675 0.7350 ;
        RECT 0.5775 0.4725 0.8925 0.5775 ;
        RECT 0.4275 0.4725 0.5025 0.7350 ;
        RECT 0.3675 0.4725 0.4275 0.5775 ;
        RECT 0.0975 0.4725 0.2925 0.6750 ;
        RECT 0.0600 0.1500 0.1500 0.3150 ;
    END
END OAI33_0011


MACRO OAI33_0111
    CLASS CORE ;
    FOREIGN OAI33_0111 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.5200 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 1.6275 0.2925 1.9425 0.7875 ;
        VIA 1.7850 0.3750 VIA12_slot ;
        VIA 1.7850 0.7050 VIA12_slot ;
        END
    END ZN
    PIN B3
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.9000 0.7125 1.3500 0.7875 ;
        RECT 0.8250 0.6825 0.9000 0.7875 ;
        VIA 0.9375 0.7500 VIA12_square ;
        END
    END B3
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.0125 0.5625 1.4775 0.6375 ;
        VIA 1.1250 0.6000 VIA12_square ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.0275 0.2625 1.4925 0.3375 ;
        VIA 1.3800 0.3000 VIA12_square ;
        END
    END B1
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.7500 0.4125 1.1775 0.4875 ;
        RECT 0.6450 0.4125 0.7500 0.6375 ;
        VIA 0.6975 0.5550 VIA12_square ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.0600 0.7125 0.5250 0.7875 ;
        VIA 0.4125 0.7500 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.0600 0.5625 0.5250 0.6375 ;
        VIA 0.2400 0.6000 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 2.2650 -0.0750 2.5200 0.0750 ;
        RECT 2.1450 -0.0750 2.2650 0.2100 ;
        RECT 1.8225 -0.0750 2.1450 0.0750 ;
        RECT 1.7475 -0.0750 1.8225 0.2325 ;
        RECT 1.4250 -0.0750 1.7475 0.0750 ;
        RECT 1.3050 -0.0750 1.4250 0.1875 ;
        RECT 1.0050 -0.0750 1.3050 0.0750 ;
        RECT 0.8850 -0.0750 1.0050 0.1875 ;
        RECT 0.0000 -0.0750 0.8850 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 2.2650 0.9750 2.5200 1.1250 ;
        RECT 2.1450 0.8625 2.2650 1.1250 ;
        RECT 1.8450 0.9750 2.1450 1.1250 ;
        RECT 1.7250 0.8550 1.8450 1.1250 ;
        RECT 1.4175 0.9750 1.7250 1.1250 ;
        RECT 1.3125 0.8325 1.4175 1.1250 ;
        RECT 0.1425 0.9750 1.3125 1.1250 ;
        RECT 0.0675 0.7950 0.1425 1.1250 ;
        RECT 0.0000 0.9750 0.0675 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 2.3850 0.2925 2.4450 0.3525 ;
        RECT 2.3850 0.8175 2.4450 0.8775 ;
        RECT 2.2725 0.4950 2.3325 0.5550 ;
        RECT 2.1750 0.1425 2.2350 0.2025 ;
        RECT 2.1750 0.8625 2.2350 0.9225 ;
        RECT 2.0700 0.4950 2.1300 0.5550 ;
        RECT 1.9650 0.2700 2.0250 0.3300 ;
        RECT 1.9650 0.7650 2.0250 0.8250 ;
        RECT 1.8600 0.4950 1.9200 0.5550 ;
        RECT 1.7550 0.1425 1.8150 0.2025 ;
        RECT 1.7550 0.8625 1.8150 0.9225 ;
        RECT 1.6500 0.4950 1.7100 0.5550 ;
        RECT 1.5450 0.2700 1.6050 0.3300 ;
        RECT 1.5450 0.7650 1.6050 0.8250 ;
        RECT 1.4400 0.4950 1.5000 0.5550 ;
        RECT 1.3350 0.1200 1.3950 0.1800 ;
        RECT 1.3350 0.8625 1.3950 0.9225 ;
        RECT 1.2375 0.4800 1.2975 0.5400 ;
        RECT 1.1250 0.1725 1.1850 0.2325 ;
        RECT 1.0200 0.4950 1.0800 0.5550 ;
        RECT 0.9150 0.1275 0.9750 0.1875 ;
        RECT 0.8175 0.4800 0.8775 0.5400 ;
        RECT 0.7050 0.1575 0.7650 0.2175 ;
        RECT 0.7050 0.8175 0.7650 0.8775 ;
        RECT 0.6000 0.4950 0.6600 0.5550 ;
        RECT 0.4950 0.3075 0.5550 0.3675 ;
        RECT 0.3900 0.4950 0.4500 0.5550 ;
        RECT 0.2850 0.1575 0.3450 0.2175 ;
        RECT 0.1800 0.4950 0.2400 0.5550 ;
        RECT 0.0750 0.2325 0.1350 0.2925 ;
        RECT 0.0750 0.8325 0.1350 0.8925 ;
        LAYER M1 ;
        RECT 2.4075 0.2850 2.4825 0.9000 ;
        RECT 2.1825 0.2850 2.4075 0.3600 ;
        RECT 2.3625 0.7950 2.4075 0.9000 ;
        RECT 2.2575 0.4650 2.3325 0.7200 ;
        RECT 2.2425 0.6450 2.2575 0.7200 ;
        RECT 2.1075 0.6450 2.2425 0.7875 ;
        RECT 2.1075 0.2850 2.1825 0.5700 ;
        RECT 1.5225 0.4950 2.1075 0.5700 ;
        RECT 1.9575 0.2175 2.0325 0.4200 ;
        RECT 1.9425 0.6675 2.0325 0.8550 ;
        RECT 1.6125 0.3300 1.9575 0.4200 ;
        RECT 1.6275 0.6675 1.9425 0.7575 ;
        RECT 1.5225 0.6675 1.6275 0.8550 ;
        RECT 1.5375 0.2175 1.6125 0.4200 ;
        RECT 1.4100 0.4950 1.5225 0.5925 ;
        RECT 1.3125 0.2625 1.4625 0.4125 ;
        RECT 1.2975 0.2625 1.3125 0.5850 ;
        RECT 1.2375 0.3375 1.2975 0.5850 ;
        RECT 1.1550 0.1500 1.2075 0.2550 ;
        RECT 1.0575 0.4650 1.1625 0.7275 ;
        RECT 1.0800 0.1500 1.1550 0.3375 ;
        RECT 0.8100 0.2625 1.0800 0.3375 ;
        RECT 0.9900 0.4650 1.0575 0.5700 ;
        RECT 0.9000 0.6450 0.9825 0.8700 ;
        RECT 0.8625 0.4500 0.9000 0.8700 ;
        RECT 0.8175 0.4500 0.8625 0.7200 ;
        RECT 0.7350 0.1500 0.8100 0.3375 ;
        RECT 0.6900 0.7950 0.7875 0.9000 ;
        RECT 0.5475 0.4500 0.7425 0.6375 ;
        RECT 0.2550 0.1500 0.7350 0.2250 ;
        RECT 0.5475 0.7125 0.6900 0.9000 ;
        RECT 0.1425 0.3000 0.6225 0.3750 ;
        RECT 0.3675 0.4725 0.4725 0.8325 ;
        RECT 0.2175 0.4500 0.2925 0.8400 ;
        RECT 0.1800 0.4500 0.2175 0.6825 ;
        RECT 0.0675 0.2025 0.1425 0.3750 ;
        LAYER VIA1 ;
        RECT 2.2575 0.5550 2.3325 0.6300 ;
        RECT 0.6600 0.8100 0.7350 0.8850 ;
        RECT 0.4425 0.3000 0.5175 0.3750 ;
        LAYER M2 ;
        RECT 2.1675 0.5550 2.3775 0.6300 ;
        RECT 2.0925 0.1125 2.1675 0.9375 ;
        RECT 0.5325 0.1125 2.0925 0.1875 ;
        RECT 0.7500 0.8625 2.0925 0.9375 ;
        RECT 0.6450 0.7725 0.7500 0.9375 ;
        RECT 0.4275 0.1125 0.5325 0.4125 ;
    END
END OAI33_0111


MACRO OAI33_1000
    CLASS CORE ;
    FOREIGN OAI33_1000 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.6800 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 0.7725 0.7125 0.8625 0.7875 ;
        RECT 0.6975 0.1125 0.7725 0.7875 ;
        RECT 0.2325 0.1125 0.6975 0.1875 ;
        VIA 0.7800 0.7500 VIA12_square ;
        VIA 0.7350 0.3375 VIA12_square ;
        END
    END ZN
    PIN B3
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.0575 0.6900 1.1625 0.9375 ;
        RECT 0.6075 0.8625 1.0575 0.9375 ;
        VIA 1.1100 0.7650 VIA12_square ;
        END
    END B3
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.2750 0.2625 1.6200 0.3375 ;
        RECT 1.1700 0.2625 1.2750 0.5775 ;
        RECT 1.0425 0.2625 1.1700 0.3375 ;
        VIA 1.2225 0.4950 VIA12_square ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.5225 0.3675 1.6275 0.6825 ;
        RECT 1.4400 0.4650 1.5225 0.5850 ;
        END
    END B1
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.9225 0.1125 1.3875 0.1875 ;
        RECT 0.9225 0.4725 0.9525 0.6375 ;
        RECT 0.8475 0.1125 0.9225 0.6375 ;
        VIA 0.9000 0.5550 VIA12_square ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.1125 0.7125 0.5775 0.7875 ;
        VIA 0.4200 0.7500 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.1125 0.5625 0.5775 0.6375 ;
        VIA 0.2400 0.6000 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.6125 -0.0750 1.6800 0.0750 ;
        RECT 1.5375 -0.0750 1.6125 0.2475 ;
        RECT 1.2150 -0.0750 1.5375 0.0750 ;
        RECT 1.0950 -0.0750 1.2150 0.1875 ;
        RECT 0.0000 -0.0750 1.0950 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.6275 0.9750 1.6800 1.1250 ;
        RECT 1.5225 0.7950 1.6275 1.1250 ;
        RECT 0.1425 0.9750 1.5225 1.1250 ;
        RECT 0.0675 0.7950 0.1425 1.1250 ;
        RECT 0.0000 0.9750 0.0675 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.5450 0.1575 1.6050 0.2175 ;
        RECT 1.5450 0.8250 1.6050 0.8850 ;
        RECT 1.4400 0.4950 1.5000 0.5550 ;
        RECT 1.3350 0.1800 1.3950 0.2400 ;
        RECT 1.2300 0.4800 1.2900 0.5400 ;
        RECT 1.1250 0.1275 1.1850 0.1875 ;
        RECT 1.0275 0.4950 1.0875 0.5550 ;
        RECT 0.9150 0.1575 0.9750 0.2175 ;
        RECT 0.9150 0.8175 0.9750 0.8775 ;
        RECT 0.7050 0.1575 0.7650 0.2175 ;
        RECT 0.7050 0.8175 0.7650 0.8775 ;
        RECT 0.6000 0.4950 0.6600 0.5550 ;
        RECT 0.4950 0.3075 0.5550 0.3675 ;
        RECT 0.3900 0.4950 0.4500 0.5550 ;
        RECT 0.2850 0.1575 0.3450 0.2175 ;
        RECT 0.1800 0.4950 0.2400 0.5550 ;
        RECT 0.0750 0.1800 0.1350 0.2400 ;
        RECT 0.0750 0.8325 0.1350 0.8925 ;
        LAYER M1 ;
        RECT 1.3125 0.1500 1.4175 0.3375 ;
        RECT 1.2225 0.4125 1.3275 0.7650 ;
        RECT 1.0200 0.2625 1.3125 0.3375 ;
        RECT 1.1850 0.4125 1.2225 0.5775 ;
        RECT 1.1100 0.6450 1.1475 0.8700 ;
        RECT 1.0725 0.4650 1.1100 0.8700 ;
        RECT 1.0275 0.4650 1.0725 0.7200 ;
        RECT 0.9450 0.1500 1.0200 0.3375 ;
        RECT 0.8625 0.7950 0.9975 0.9000 ;
        RECT 0.8475 0.4725 0.9525 0.6375 ;
        RECT 0.2550 0.1500 0.9450 0.2250 ;
        RECT 0.6600 0.7125 0.8625 0.9000 ;
        RECT 0.5700 0.4725 0.8475 0.5925 ;
        RECT 0.1500 0.3000 0.8175 0.3750 ;
        RECT 0.3675 0.4725 0.4725 0.8325 ;
        RECT 0.2175 0.4500 0.2925 0.8400 ;
        RECT 0.1800 0.4500 0.2175 0.6825 ;
        RECT 0.0450 0.1500 0.1500 0.3750 ;
    END
END OAI33_1000


MACRO OAI33_1010
    CLASS CORE ;
    FOREIGN OAI33_1010 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.6800 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 0.7725 0.7125 0.8625 0.7875 ;
        RECT 0.6975 0.1125 0.7725 0.7875 ;
        RECT 0.2325 0.1125 0.6975 0.1875 ;
        VIA 0.7800 0.7500 VIA12_square ;
        VIA 0.7350 0.3375 VIA12_square ;
        END
    END ZN
    PIN B3
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.0575 0.6900 1.1625 0.9375 ;
        RECT 0.6075 0.8625 1.0575 0.9375 ;
        VIA 1.1100 0.7650 VIA12_square ;
        END
    END B3
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.2750 0.2625 1.6200 0.3375 ;
        RECT 1.1700 0.2625 1.2750 0.5775 ;
        RECT 1.0425 0.2625 1.1700 0.3375 ;
        VIA 1.2225 0.4950 VIA12_square ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.5225 0.3675 1.6275 0.6825 ;
        RECT 1.4400 0.4650 1.5225 0.5850 ;
        END
    END B1
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.9225 0.1125 1.3875 0.1875 ;
        RECT 0.9225 0.4725 0.9525 0.6375 ;
        RECT 0.8475 0.1125 0.9225 0.6375 ;
        VIA 0.9000 0.5550 VIA12_square ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.1125 0.7125 0.5775 0.7875 ;
        VIA 0.4200 0.7500 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.1125 0.5625 0.5775 0.6375 ;
        VIA 0.2400 0.6000 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.6125 -0.0750 1.6800 0.0750 ;
        RECT 1.5375 -0.0750 1.6125 0.2475 ;
        RECT 1.2150 -0.0750 1.5375 0.0750 ;
        RECT 1.0950 -0.0750 1.2150 0.1875 ;
        RECT 0.0000 -0.0750 1.0950 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.6275 0.9750 1.6800 1.1250 ;
        RECT 1.5225 0.7950 1.6275 1.1250 ;
        RECT 0.1425 0.9750 1.5225 1.1250 ;
        RECT 0.0675 0.7950 0.1425 1.1250 ;
        RECT 0.0000 0.9750 0.0675 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.5450 0.1575 1.6050 0.2175 ;
        RECT 1.5450 0.8250 1.6050 0.8850 ;
        RECT 1.4400 0.4950 1.5000 0.5550 ;
        RECT 1.3350 0.1800 1.3950 0.2400 ;
        RECT 1.2300 0.4800 1.2900 0.5400 ;
        RECT 1.1250 0.1275 1.1850 0.1875 ;
        RECT 1.0275 0.4950 1.0875 0.5550 ;
        RECT 0.9150 0.1575 0.9750 0.2175 ;
        RECT 0.9150 0.8175 0.9750 0.8775 ;
        RECT 0.7050 0.1575 0.7650 0.2175 ;
        RECT 0.7050 0.8175 0.7650 0.8775 ;
        RECT 0.6000 0.4950 0.6600 0.5550 ;
        RECT 0.4950 0.3075 0.5550 0.3675 ;
        RECT 0.3900 0.4950 0.4500 0.5550 ;
        RECT 0.2850 0.1575 0.3450 0.2175 ;
        RECT 0.1800 0.4950 0.2400 0.5550 ;
        RECT 0.0750 0.1800 0.1350 0.2400 ;
        RECT 0.0750 0.8325 0.1350 0.8925 ;
        LAYER M1 ;
        RECT 1.3125 0.1500 1.4175 0.3375 ;
        RECT 1.2225 0.4125 1.3275 0.7650 ;
        RECT 1.0200 0.2625 1.3125 0.3375 ;
        RECT 1.1850 0.4125 1.2225 0.5775 ;
        RECT 1.1100 0.6450 1.1475 0.8700 ;
        RECT 1.0725 0.4650 1.1100 0.8700 ;
        RECT 1.0275 0.4650 1.0725 0.7200 ;
        RECT 0.9450 0.1500 1.0200 0.3375 ;
        RECT 0.8625 0.7950 0.9975 0.9000 ;
        RECT 0.8475 0.4725 0.9525 0.6375 ;
        RECT 0.2550 0.1500 0.9450 0.2250 ;
        RECT 0.6600 0.7125 0.8625 0.9000 ;
        RECT 0.5700 0.4725 0.8475 0.5925 ;
        RECT 0.1500 0.3000 0.8175 0.3750 ;
        RECT 0.3675 0.4725 0.4725 0.8325 ;
        RECT 0.2175 0.4500 0.2925 0.8400 ;
        RECT 0.1800 0.4500 0.2175 0.6825 ;
        RECT 0.0450 0.1500 0.1500 0.3750 ;
    END
END OAI33_1010


MACRO OR2_0010
    CLASS CORE ;
    FOREIGN OR2_0010 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.2000 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 3.4125 0.2775 3.5700 0.3975 ;
        RECT 3.4125 0.6525 3.5700 0.7725 ;
        RECT 3.0975 0.2775 3.4125 0.7725 ;
        RECT 2.9400 0.2775 3.0975 0.3975 ;
        RECT 2.9400 0.6525 3.0975 0.7725 ;
        VIA 3.4125 0.3375 VIA12_slot ;
        VIA 3.4125 0.7125 VIA12_slot ;
        VIA 3.0975 0.3375 VIA12_slot ;
        VIA 3.0975 0.7125 VIA12_slot ;
        END
    END Z
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.3375 0.4575 1.3200 0.5700 ;
        RECT 0.1725 0.4125 0.3375 0.6375 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.9275 0.4125 2.0325 0.6075 ;
        RECT 1.4100 0.4125 1.9275 0.4875 ;
        VIA 1.9800 0.5100 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 4.1550 -0.0750 4.2000 0.0750 ;
        RECT 4.0350 -0.0750 4.1550 0.2925 ;
        RECT 3.7350 -0.0750 4.0350 0.0750 ;
        RECT 3.6150 -0.0750 3.7350 0.2025 ;
        RECT 3.3150 -0.0750 3.6150 0.0750 ;
        RECT 3.1950 -0.0750 3.3150 0.2025 ;
        RECT 2.8950 -0.0750 3.1950 0.0750 ;
        RECT 2.7750 -0.0750 2.8950 0.2025 ;
        RECT 2.4750 -0.0750 2.7750 0.0750 ;
        RECT 2.3550 -0.0750 2.4750 0.2250 ;
        RECT 2.2650 -0.0750 2.3550 0.0750 ;
        RECT 2.1450 -0.0750 2.2650 0.2250 ;
        RECT 1.8375 -0.0750 2.1450 0.0750 ;
        RECT 1.7325 -0.0750 1.8375 0.2250 ;
        RECT 1.4175 -0.0750 1.7325 0.0750 ;
        RECT 1.3125 -0.0750 1.4175 0.2250 ;
        RECT 0.9975 -0.0750 1.3125 0.0750 ;
        RECT 0.8925 -0.0750 0.9975 0.2250 ;
        RECT 0.5850 -0.0750 0.8925 0.0750 ;
        RECT 0.4650 -0.0750 0.5850 0.1875 ;
        RECT 0.1425 -0.0750 0.4650 0.0750 ;
        RECT 0.0675 -0.0750 0.1425 0.2700 ;
        RECT 0.0000 -0.0750 0.0675 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 4.1550 0.9750 4.2000 1.1250 ;
        RECT 4.0350 0.6600 4.1550 1.1250 ;
        RECT 3.7350 0.9750 4.0350 1.1250 ;
        RECT 3.6150 0.8475 3.7350 1.1250 ;
        RECT 3.3150 0.9750 3.6150 1.1250 ;
        RECT 3.1950 0.8475 3.3150 1.1250 ;
        RECT 2.8950 0.9750 3.1950 1.1250 ;
        RECT 2.7750 0.8475 2.8950 1.1250 ;
        RECT 2.4675 0.9750 2.7750 1.1250 ;
        RECT 2.3625 0.8025 2.4675 1.1250 ;
        RECT 1.2150 0.9750 2.3625 1.1250 ;
        RECT 1.0950 0.8625 1.2150 1.1250 ;
        RECT 0.7950 0.9750 1.0950 1.1250 ;
        RECT 0.6750 0.8625 0.7950 1.1250 ;
        RECT 0.3750 0.9750 0.6750 1.1250 ;
        RECT 0.2550 0.8625 0.3750 1.1250 ;
        RECT 0.0000 0.9750 0.2550 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 4.0650 0.2175 4.1250 0.2775 ;
        RECT 4.0650 0.6675 4.1250 0.7275 ;
        RECT 4.0650 0.8325 4.1250 0.8925 ;
        RECT 3.9600 0.4800 4.0200 0.5400 ;
        RECT 3.8550 0.3075 3.9150 0.3675 ;
        RECT 3.8550 0.6825 3.9150 0.7425 ;
        RECT 3.7500 0.4800 3.8100 0.5400 ;
        RECT 3.6450 0.1350 3.7050 0.1950 ;
        RECT 3.6450 0.8550 3.7050 0.9150 ;
        RECT 3.5400 0.4800 3.6000 0.5400 ;
        RECT 3.4350 0.3075 3.4950 0.3675 ;
        RECT 3.4350 0.6825 3.4950 0.7425 ;
        RECT 3.3300 0.4800 3.3900 0.5400 ;
        RECT 3.2250 0.1350 3.2850 0.1950 ;
        RECT 3.2250 0.8550 3.2850 0.9150 ;
        RECT 3.1200 0.4800 3.1800 0.5400 ;
        RECT 3.0150 0.3075 3.0750 0.3675 ;
        RECT 3.0150 0.6825 3.0750 0.7425 ;
        RECT 2.9100 0.4800 2.9700 0.5400 ;
        RECT 2.8050 0.1350 2.8650 0.1950 ;
        RECT 2.8050 0.8550 2.8650 0.9150 ;
        RECT 2.7000 0.4800 2.7600 0.5400 ;
        RECT 2.5950 0.3075 2.6550 0.3675 ;
        RECT 2.5950 0.6825 2.6550 0.7425 ;
        RECT 2.4900 0.4800 2.5500 0.5400 ;
        RECT 2.3850 0.1575 2.4450 0.2175 ;
        RECT 2.3850 0.8325 2.4450 0.8925 ;
        RECT 2.1750 0.1575 2.2350 0.2175 ;
        RECT 2.1750 0.8175 2.2350 0.8775 ;
        RECT 2.0700 0.4800 2.1300 0.5400 ;
        RECT 1.9650 0.2100 2.0250 0.2700 ;
        RECT 1.9650 0.6750 2.0250 0.7350 ;
        RECT 1.8600 0.4800 1.9200 0.5400 ;
        RECT 1.7550 0.1350 1.8150 0.1950 ;
        RECT 1.7550 0.8325 1.8150 0.8925 ;
        RECT 1.6500 0.4800 1.7100 0.5400 ;
        RECT 1.5450 0.3075 1.6050 0.3675 ;
        RECT 1.5450 0.6750 1.6050 0.7350 ;
        RECT 1.4400 0.4800 1.5000 0.5400 ;
        RECT 1.3350 0.1350 1.3950 0.1950 ;
        RECT 1.3350 0.8325 1.3950 0.8925 ;
        RECT 1.2300 0.4800 1.2900 0.5400 ;
        RECT 1.1250 0.3075 1.1850 0.3675 ;
        RECT 1.1250 0.8625 1.1850 0.9225 ;
        RECT 1.0200 0.4800 1.0800 0.5400 ;
        RECT 0.9150 0.1350 0.9750 0.1950 ;
        RECT 0.9150 0.7200 0.9750 0.7800 ;
        RECT 0.8100 0.4800 0.8700 0.5400 ;
        RECT 0.7050 0.1800 0.7650 0.2400 ;
        RECT 0.7050 0.8625 0.7650 0.9225 ;
        RECT 0.6000 0.4800 0.6600 0.5400 ;
        RECT 0.4950 0.1275 0.5550 0.1875 ;
        RECT 0.4950 0.7200 0.5550 0.7800 ;
        RECT 0.3900 0.4800 0.4500 0.5400 ;
        RECT 0.0750 0.7800 0.1350 0.8400 ;
        RECT 0.2850 0.1800 0.3450 0.2400 ;
        RECT 0.2850 0.8625 0.3450 0.9225 ;
        RECT 0.1800 0.4800 0.2400 0.5400 ;
        RECT 0.0750 0.1575 0.1350 0.2175 ;
        LAYER M1 ;
        RECT 2.4525 0.4725 4.0950 0.5475 ;
        RECT 2.5875 0.2775 3.9300 0.3975 ;
        RECT 2.5875 0.6525 3.9300 0.7725 ;
        RECT 2.3775 0.3000 2.4525 0.7200 ;
        RECT 2.0325 0.3000 2.3775 0.3750 ;
        RECT 2.0550 0.6450 2.3775 0.7200 ;
        RECT 2.1525 0.7950 2.2575 0.9000 ;
        RECT 1.4100 0.4575 2.1975 0.5700 ;
        RECT 1.3650 0.8250 2.1525 0.9000 ;
        RECT 1.5150 0.6450 2.0550 0.7500 ;
        RECT 1.9575 0.1800 2.0325 0.3750 ;
        RECT 0.7875 0.3000 1.9575 0.3750 ;
        RECT 1.2900 0.7125 1.3650 0.9000 ;
        RECT 0.1425 0.7125 1.2900 0.7875 ;
        RECT 0.6825 0.1500 0.7875 0.3750 ;
        RECT 0.3675 0.2625 0.6825 0.3375 ;
        RECT 0.2625 0.1500 0.3675 0.3375 ;
        RECT 0.0675 0.7125 0.1425 0.8700 ;
        LAYER M2 ;
        RECT 3.4425 0.2775 3.5700 0.3975 ;
        RECT 3.4425 0.6525 3.5700 0.7725 ;
        RECT 2.9400 0.2775 3.0675 0.3975 ;
        RECT 2.9400 0.6525 3.0675 0.7725 ;
    END
END OR2_0010


MACRO OR2_0011
    CLASS CORE ;
    FOREIGN OR2_0011 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.0500 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.9375 0.3075 1.0125 0.7350 ;
        RECT 0.7725 0.3075 0.9375 0.3825 ;
        RECT 0.7725 0.6600 0.9375 0.7350 ;
        RECT 0.6975 0.2175 0.7725 0.3825 ;
        RECT 0.6975 0.6600 0.7725 0.8325 ;
        END
    END Z
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.4500 0.1125 0.9150 0.1875 ;
        RECT 0.4500 0.4050 0.4800 0.5700 ;
        RECT 0.3750 0.1125 0.4500 0.5700 ;
        VIA 0.4275 0.4875 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1425 0.4500 0.2325 0.5700 ;
        RECT 0.0675 0.3675 0.1425 0.6825 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.0050 -0.0750 1.0500 0.0750 ;
        RECT 0.8850 -0.0750 1.0050 0.2325 ;
        RECT 0.5850 -0.0750 0.8850 0.0750 ;
        RECT 0.4650 -0.0750 0.5850 0.1800 ;
        RECT 0.1500 -0.0750 0.4650 0.0750 ;
        RECT 0.0675 -0.0750 0.1500 0.2475 ;
        RECT 0.0000 -0.0750 0.0675 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.9975 0.9750 1.0500 1.1250 ;
        RECT 0.8925 0.8100 0.9975 1.1250 ;
        RECT 0.5850 0.9750 0.8925 1.1250 ;
        RECT 0.4650 0.8700 0.5850 1.1250 ;
        RECT 0.0000 0.9750 0.4650 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 0.9150 0.1650 0.9750 0.2250 ;
        RECT 0.9150 0.8325 0.9750 0.8925 ;
        RECT 0.8025 0.4875 0.8625 0.5475 ;
        RECT 0.7050 0.2700 0.7650 0.3300 ;
        RECT 0.7050 0.7200 0.7650 0.7800 ;
        RECT 0.6000 0.4875 0.6600 0.5475 ;
        RECT 0.4950 0.1200 0.5550 0.1800 ;
        RECT 0.4950 0.8700 0.5550 0.9300 ;
        RECT 0.3900 0.4875 0.4500 0.5475 ;
        RECT 0.2850 0.1800 0.3450 0.2400 ;
        RECT 0.1725 0.4800 0.2325 0.5400 ;
        RECT 0.0750 0.1575 0.1350 0.2175 ;
        RECT 0.0750 0.8175 0.1350 0.8775 ;
        LAYER M1 ;
        RECT 0.6225 0.4575 0.8625 0.5775 ;
        RECT 0.5475 0.2550 0.6225 0.7950 ;
        RECT 0.3675 0.2550 0.5475 0.3300 ;
        RECT 0.3900 0.7200 0.5475 0.7950 ;
        RECT 0.3075 0.4050 0.4725 0.6450 ;
        RECT 0.3150 0.7200 0.3900 0.9000 ;
        RECT 0.2625 0.1575 0.3675 0.3300 ;
        RECT 0.0525 0.7950 0.3150 0.9000 ;
    END
END OR2_0011


MACRO OR2_0100
    CLASS CORE ;
    FOREIGN OR2_0100 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.1500 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 2.3625 0.2625 2.5200 0.3825 ;
        RECT 2.3625 0.6600 2.5200 0.7800 ;
        RECT 2.0475 0.2625 2.3625 0.7800 ;
        RECT 1.8900 0.2625 2.0475 0.3825 ;
        RECT 1.8900 0.6600 2.0475 0.7800 ;
        VIA 2.3625 0.3225 VIA12_slot ;
        VIA 2.3625 0.7200 VIA12_slot ;
        VIA 2.0475 0.3225 VIA12_slot ;
        VIA 2.0475 0.7200 VIA12_slot ;
        END
    END Z
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.2000 0.2625 1.2750 0.5850 ;
        RECT 0.7350 0.2625 1.2000 0.3375 ;
        RECT 0.6600 0.2625 0.7350 0.5550 ;
        RECT 0.5775 0.4500 0.6600 0.5550 ;
        VIA 1.2375 0.5025 VIA12_square ;
        VIA 0.6525 0.5025 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.9450 0.4575 1.0200 0.5625 ;
        RECT 0.8700 0.4575 0.9450 0.7875 ;
        RECT 0.5025 0.7125 0.8700 0.7875 ;
        RECT 0.4275 0.5625 0.5025 0.7875 ;
        RECT 0.0975 0.5625 0.4275 0.6375 ;
        VIA 0.9450 0.5100 VIA12_square ;
        VIA 0.2100 0.6000 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 3.0825 -0.0750 3.1500 0.0750 ;
        RECT 3.0075 -0.0750 3.0825 0.2925 ;
        RECT 2.6850 -0.0750 3.0075 0.0750 ;
        RECT 2.5650 -0.0750 2.6850 0.1875 ;
        RECT 2.2650 -0.0750 2.5650 0.0750 ;
        RECT 2.1450 -0.0750 2.2650 0.1875 ;
        RECT 1.8450 -0.0750 2.1450 0.0750 ;
        RECT 1.7250 -0.0750 1.8450 0.1875 ;
        RECT 1.4250 -0.0750 1.7250 0.0750 ;
        RECT 1.3050 -0.0750 1.4250 0.1950 ;
        RECT 1.0050 -0.0750 1.3050 0.0750 ;
        RECT 0.8850 -0.0750 1.0050 0.1950 ;
        RECT 0.5850 -0.0750 0.8850 0.0750 ;
        RECT 0.4650 -0.0750 0.5850 0.1950 ;
        RECT 0.1425 -0.0750 0.4650 0.0750 ;
        RECT 0.0675 -0.0750 0.1425 0.2625 ;
        RECT 0.0000 -0.0750 0.0675 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 3.0825 0.9750 3.1500 1.1250 ;
        RECT 3.0075 0.6375 3.0825 1.1250 ;
        RECT 2.6850 0.9750 3.0075 1.1250 ;
        RECT 2.5650 0.8550 2.6850 1.1250 ;
        RECT 2.2650 0.9750 2.5650 1.1250 ;
        RECT 2.1450 0.8550 2.2650 1.1250 ;
        RECT 1.8450 0.9750 2.1450 1.1250 ;
        RECT 1.7250 0.8550 1.8450 1.1250 ;
        RECT 1.4250 0.9750 1.7250 1.1250 ;
        RECT 1.3050 0.8625 1.4250 1.1250 ;
        RECT 0.5850 0.9750 1.3050 1.1250 ;
        RECT 0.4650 0.8625 0.5850 1.1250 ;
        RECT 0.0000 0.9750 0.4650 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 3.0150 0.1875 3.0750 0.2475 ;
        RECT 3.0150 0.6675 3.0750 0.7275 ;
        RECT 3.0150 0.8325 3.0750 0.8925 ;
        RECT 2.9100 0.4650 2.9700 0.5250 ;
        RECT 2.8050 0.2850 2.8650 0.3450 ;
        RECT 2.8050 0.6900 2.8650 0.7500 ;
        RECT 2.7000 0.4650 2.7600 0.5250 ;
        RECT 2.5950 0.1275 2.6550 0.1875 ;
        RECT 2.5950 0.8625 2.6550 0.9225 ;
        RECT 2.4900 0.4650 2.5500 0.5250 ;
        RECT 2.3850 0.2850 2.4450 0.3450 ;
        RECT 2.3850 0.6900 2.4450 0.7500 ;
        RECT 2.2800 0.4650 2.3400 0.5250 ;
        RECT 2.1750 0.1275 2.2350 0.1875 ;
        RECT 2.1750 0.8625 2.2350 0.9225 ;
        RECT 2.0700 0.4650 2.1300 0.5250 ;
        RECT 1.9650 0.2850 2.0250 0.3450 ;
        RECT 1.9650 0.6900 2.0250 0.7500 ;
        RECT 1.8600 0.4650 1.9200 0.5250 ;
        RECT 1.7550 0.1275 1.8150 0.1875 ;
        RECT 1.7550 0.8625 1.8150 0.9225 ;
        RECT 1.6500 0.4650 1.7100 0.5250 ;
        RECT 1.5450 0.2925 1.6050 0.3525 ;
        RECT 1.5450 0.6900 1.6050 0.7500 ;
        RECT 1.4400 0.4650 1.5000 0.5250 ;
        RECT 1.3350 0.1275 1.3950 0.1875 ;
        RECT 1.3350 0.8625 1.3950 0.9225 ;
        RECT 1.2300 0.4800 1.2900 0.5400 ;
        RECT 1.1250 0.1725 1.1850 0.2325 ;
        RECT 1.0200 0.4650 1.0800 0.5250 ;
        RECT 0.9150 0.1275 0.9750 0.1875 ;
        RECT 0.9150 0.7200 0.9750 0.7800 ;
        RECT 0.8100 0.4650 0.8700 0.5250 ;
        RECT 0.7050 0.1725 0.7650 0.2325 ;
        RECT 0.6000 0.4650 0.6600 0.5250 ;
        RECT 0.4950 0.1275 0.5550 0.1875 ;
        RECT 0.4950 0.8625 0.5550 0.9225 ;
        RECT 0.3900 0.4650 0.4500 0.5250 ;
        RECT 0.2850 0.1725 0.3450 0.2325 ;
        RECT 0.1800 0.4650 0.2400 0.5250 ;
        RECT 0.0750 0.1575 0.1350 0.2175 ;
        RECT 0.0750 0.7425 0.1350 0.8025 ;
        LAYER M1 ;
        RECT 1.4625 0.4575 3.0000 0.5325 ;
        RECT 1.5375 0.2625 2.8875 0.3825 ;
        RECT 1.5375 0.6600 2.8875 0.7800 ;
        RECT 1.3875 0.2700 1.4625 0.7875 ;
        RECT 1.2150 0.2700 1.3875 0.3450 ;
        RECT 0.1425 0.7125 1.3875 0.7875 ;
        RECT 1.1625 0.4200 1.3125 0.6300 ;
        RECT 1.0950 0.1500 1.2150 0.3450 ;
        RECT 0.7875 0.2700 1.0950 0.3450 ;
        RECT 0.8025 0.4350 1.0875 0.6075 ;
        RECT 0.6825 0.1500 0.7875 0.3450 ;
        RECT 0.3825 0.4350 0.7275 0.5550 ;
        RECT 0.3675 0.2700 0.6825 0.3450 ;
        RECT 0.2625 0.1500 0.3675 0.3450 ;
        RECT 0.1275 0.4200 0.2925 0.6375 ;
        RECT 0.0675 0.7125 0.1425 0.8325 ;
        LAYER M2 ;
        RECT 2.3925 0.2625 2.5200 0.3825 ;
        RECT 2.3925 0.6600 2.5200 0.7800 ;
        RECT 1.8900 0.2625 2.0175 0.3825 ;
        RECT 1.8900 0.6600 2.0175 0.7800 ;
    END
END OR2_0100


MACRO OR2_0111
    CLASS CORE ;
    FOREIGN OR2_0111 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.8900 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 1.2075 0.2400 1.5225 0.7500 ;
        VIA 1.3650 0.3225 VIA12_slot ;
        VIA 1.3650 0.6675 VIA12_slot ;
        END
    END Z
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.8025 0.2625 0.9075 0.6075 ;
        RECT 0.3525 0.2625 0.8025 0.3375 ;
        RECT 0.2775 0.2625 0.3525 0.4875 ;
        RECT 0.1125 0.4125 0.2775 0.4875 ;
        VIA 0.8550 0.5250 VIA12_square ;
        VIA 0.2250 0.4500 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.5925 0.7125 1.0575 0.7875 ;
        RECT 0.4875 0.4275 0.5925 0.7875 ;
        VIA 0.5400 0.5025 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.8225 -0.0750 1.8900 0.0750 ;
        RECT 1.7475 -0.0750 1.8225 0.3150 ;
        RECT 1.4250 -0.0750 1.7475 0.0750 ;
        RECT 1.3050 -0.0750 1.4250 0.1950 ;
        RECT 1.0050 -0.0750 1.3050 0.0750 ;
        RECT 0.8850 -0.0750 1.0050 0.1875 ;
        RECT 0.5850 -0.0750 0.8850 0.0750 ;
        RECT 0.4650 -0.0750 0.5850 0.1875 ;
        RECT 0.1575 -0.0750 0.4650 0.0750 ;
        RECT 0.0525 -0.0750 0.1575 0.2625 ;
        RECT 0.0000 -0.0750 0.0525 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.8225 0.9750 1.8900 1.1250 ;
        RECT 1.7475 0.6375 1.8225 1.1250 ;
        RECT 1.4025 0.9750 1.7475 1.1250 ;
        RECT 1.3275 0.8175 1.4025 1.1250 ;
        RECT 1.0050 0.9750 1.3275 1.1250 ;
        RECT 0.8850 0.8550 1.0050 1.1250 ;
        RECT 0.1575 0.9750 0.8850 1.1250 ;
        RECT 0.0525 0.6450 0.1575 1.1250 ;
        RECT 0.0000 0.9750 0.0525 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.7550 0.2250 1.8150 0.2850 ;
        RECT 1.7550 0.6675 1.8150 0.7275 ;
        RECT 1.7550 0.8325 1.8150 0.8925 ;
        RECT 1.6500 0.4650 1.7100 0.5250 ;
        RECT 1.5450 0.2250 1.6050 0.2850 ;
        RECT 1.5450 0.7575 1.6050 0.8175 ;
        RECT 1.4400 0.4650 1.5000 0.5250 ;
        RECT 1.3350 0.1275 1.3950 0.1875 ;
        RECT 1.3350 0.8475 1.3950 0.9075 ;
        RECT 1.2300 0.4650 1.2900 0.5250 ;
        RECT 1.1250 0.2250 1.1850 0.2850 ;
        RECT 1.1250 0.7575 1.1850 0.8175 ;
        RECT 1.0200 0.4650 1.0800 0.5250 ;
        RECT 0.9150 0.1275 0.9750 0.1875 ;
        RECT 0.9150 0.8625 0.9750 0.9225 ;
        RECT 0.8100 0.4800 0.8700 0.5400 ;
        RECT 0.7050 0.1725 0.7650 0.2325 ;
        RECT 0.6000 0.4650 0.6600 0.5250 ;
        RECT 0.4950 0.1275 0.5550 0.1875 ;
        RECT 0.4950 0.7125 0.5550 0.7725 ;
        RECT 0.3900 0.4650 0.4500 0.5250 ;
        RECT 0.2850 0.1725 0.3450 0.2325 ;
        RECT 0.1800 0.4650 0.2400 0.5250 ;
        RECT 0.0750 0.1575 0.1350 0.2175 ;
        RECT 0.0750 0.6675 0.1350 0.7275 ;
        RECT 0.0750 0.8325 0.1350 0.8925 ;
        LAYER M1 ;
        RECT 1.0425 0.4425 1.7400 0.5475 ;
        RECT 1.5225 0.1950 1.6275 0.3675 ;
        RECT 1.5375 0.6225 1.6125 0.8700 ;
        RECT 1.1925 0.6225 1.5375 0.7125 ;
        RECT 1.2075 0.2775 1.5225 0.3675 ;
        RECT 1.1175 0.1950 1.2075 0.3675 ;
        RECT 1.1175 0.6225 1.1925 0.8700 ;
        RECT 0.9675 0.2625 1.0425 0.7800 ;
        RECT 0.7950 0.2625 0.9675 0.3375 ;
        RECT 0.4575 0.7050 0.9675 0.7800 ;
        RECT 0.7425 0.4200 0.8925 0.6300 ;
        RECT 0.6750 0.1500 0.7950 0.3375 ;
        RECT 0.3750 0.2625 0.6750 0.3375 ;
        RECT 0.3825 0.4350 0.6675 0.5625 ;
        RECT 0.2550 0.1500 0.3750 0.3375 ;
        RECT 0.0750 0.4125 0.3075 0.5700 ;
    END
END OR2_0111


MACRO OR2_1000
    CLASS CORE ;
    FOREIGN OR2_1000 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.8400 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1425 0.1500 0.1650 0.2250 ;
        RECT 0.1125 0.6675 0.1575 0.9000 ;
        RECT 0.1125 0.1500 0.1425 0.3825 ;
        RECT 0.0375 0.1500 0.1125 0.9000 ;
        END
    END Z
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.1875 0.5625 0.6825 0.6375 ;
        VIA 0.4050 0.6000 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.4575 0.7125 0.7725 0.7875 ;
        RECT 0.3825 0.7125 0.4575 0.9375 ;
        RECT 0.0675 0.8625 0.3825 0.9375 ;
        VIA 0.5700 0.7500 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.8025 -0.0750 0.8400 0.0750 ;
        RECT 0.6600 -0.0750 0.8025 0.2250 ;
        RECT 0.3750 -0.0750 0.6600 0.0750 ;
        RECT 0.2700 -0.0750 0.3750 0.2250 ;
        RECT 0.0000 -0.0750 0.2700 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.3750 0.9750 0.8400 1.1250 ;
        RECT 0.2550 0.8400 0.3750 1.1250 ;
        RECT 0.0000 0.9750 0.2550 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 0.7050 0.1575 0.7650 0.2175 ;
        RECT 0.7050 0.8175 0.7650 0.8775 ;
        RECT 0.5925 0.4950 0.6525 0.5550 ;
        RECT 0.4950 0.1725 0.5550 0.2325 ;
        RECT 0.3900 0.5550 0.4500 0.6150 ;
        RECT 0.2850 0.1350 0.3450 0.1950 ;
        RECT 0.2850 0.8550 0.3450 0.9150 ;
        RECT 0.1875 0.4800 0.2475 0.5400 ;
        RECT 0.0750 0.1575 0.1350 0.2175 ;
        RECT 0.0750 0.8175 0.1350 0.8775 ;
        LAYER M1 ;
        RECT 0.7275 0.3000 0.8025 0.9000 ;
        RECT 0.5775 0.3000 0.7275 0.3750 ;
        RECT 0.6825 0.7950 0.7275 0.9000 ;
        RECT 0.6075 0.4500 0.6525 0.6000 ;
        RECT 0.5325 0.4500 0.6075 0.8700 ;
        RECT 0.4725 0.1500 0.5775 0.3750 ;
        RECT 0.2925 0.3000 0.4725 0.3750 ;
        RECT 0.3675 0.4800 0.4575 0.7650 ;
        RECT 0.2700 0.6900 0.3675 0.7650 ;
        RECT 0.2175 0.3000 0.2925 0.5700 ;
        RECT 0.1875 0.4500 0.2175 0.5700 ;
    END
END OR2_1000


MACRO OR2_1010
    CLASS CORE ;
    FOREIGN OR2_1010 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.8400 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1125 0.2175 0.1425 0.3825 ;
        RECT 0.1125 0.6675 0.1425 0.8325 ;
        RECT 0.0375 0.2175 0.1125 0.8325 ;
        END
    END Z
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.3675 0.4650 0.4725 0.7875 ;
        RECT 0.3075 0.7125 0.3675 0.7875 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.6225 0.4500 0.6525 0.6000 ;
        RECT 0.5475 0.4500 0.6225 0.8325 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.8025 -0.0750 0.8400 0.0750 ;
        RECT 0.6600 -0.0750 0.8025 0.2250 ;
        RECT 0.3750 -0.0750 0.6600 0.0750 ;
        RECT 0.2550 -0.0750 0.3750 0.2175 ;
        RECT 0.0000 -0.0750 0.2550 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.3750 0.9750 0.8400 1.1250 ;
        RECT 0.2550 0.8625 0.3750 1.1250 ;
        RECT 0.0000 0.9750 0.2550 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 0.7050 0.1575 0.7650 0.2175 ;
        RECT 0.7050 0.7200 0.7650 0.7800 ;
        RECT 0.5925 0.4950 0.6525 0.5550 ;
        RECT 0.4950 0.1725 0.5550 0.2325 ;
        RECT 0.3900 0.4950 0.4500 0.5550 ;
        RECT 0.2850 0.1575 0.3450 0.2175 ;
        RECT 0.2850 0.8625 0.3450 0.9225 ;
        RECT 0.1875 0.4800 0.2475 0.5400 ;
        RECT 0.0750 0.2700 0.1350 0.3300 ;
        RECT 0.0750 0.7200 0.1350 0.7800 ;
        LAYER M1 ;
        RECT 0.7275 0.3000 0.8025 0.8325 ;
        RECT 0.5775 0.3000 0.7275 0.3750 ;
        RECT 0.6975 0.6675 0.7275 0.8325 ;
        RECT 0.4725 0.1500 0.5775 0.3750 ;
        RECT 0.2925 0.3000 0.4725 0.3750 ;
        RECT 0.2175 0.3000 0.2925 0.5700 ;
        RECT 0.1875 0.4500 0.2175 0.5700 ;
    END
END OR2_1010


MACRO OR3_0011
    CLASS CORE ;
    FOREIGN OR3_0011 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.2600 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 1.1475 0.3075 1.2225 0.7350 ;
        RECT 0.9825 0.3075 1.1475 0.3825 ;
        RECT 0.9825 0.6600 1.1475 0.7350 ;
        RECT 0.9075 0.2175 0.9825 0.3825 ;
        RECT 0.9075 0.6600 0.9825 0.8325 ;
        END
    END Z
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.0675 0.4050 0.2400 0.6900 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.4575 0.7125 0.9225 0.7875 ;
        RECT 0.3825 0.3975 0.4575 0.7875 ;
        VIA 0.4200 0.5100 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.6600 0.1125 1.1250 0.1875 ;
        RECT 0.5850 0.1125 0.6600 0.5700 ;
        VIA 0.6225 0.4875 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.2150 -0.0750 1.2600 0.0750 ;
        RECT 1.0950 -0.0750 1.2150 0.2325 ;
        RECT 0.7950 -0.0750 1.0950 0.0750 ;
        RECT 0.6750 -0.0750 0.7950 0.1800 ;
        RECT 0.3750 -0.0750 0.6750 0.0750 ;
        RECT 0.2550 -0.0750 0.3750 0.1800 ;
        RECT 0.0000 -0.0750 0.2550 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.2075 0.9750 1.2600 1.1250 ;
        RECT 1.1025 0.8100 1.2075 1.1250 ;
        RECT 0.7950 0.9750 1.1025 1.1250 ;
        RECT 0.6750 0.8700 0.7950 1.1250 ;
        RECT 0.0000 0.9750 0.6750 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.1250 0.1650 1.1850 0.2250 ;
        RECT 1.1250 0.8325 1.1850 0.8925 ;
        RECT 1.0125 0.4875 1.0725 0.5475 ;
        RECT 0.9150 0.2700 0.9750 0.3300 ;
        RECT 0.9150 0.7200 0.9750 0.7800 ;
        RECT 0.8100 0.4875 0.8700 0.5475 ;
        RECT 0.7050 0.1200 0.7650 0.1800 ;
        RECT 0.7050 0.8700 0.7650 0.9300 ;
        RECT 0.6000 0.4875 0.6600 0.5475 ;
        RECT 0.4950 0.1800 0.5550 0.2400 ;
        RECT 0.3900 0.4875 0.4500 0.5475 ;
        RECT 0.2850 0.1200 0.3450 0.1800 ;
        RECT 0.1800 0.4950 0.2400 0.5550 ;
        RECT 0.0750 0.1575 0.1350 0.2175 ;
        RECT 0.0750 0.8175 0.1350 0.8775 ;
        LAYER M1 ;
        RECT 0.8325 0.4575 1.0725 0.5775 ;
        RECT 0.7575 0.2550 0.8325 0.7950 ;
        RECT 0.5775 0.2550 0.7575 0.3300 ;
        RECT 0.6000 0.7200 0.7575 0.7950 ;
        RECT 0.5400 0.4050 0.6825 0.6450 ;
        RECT 0.0450 0.7950 0.5250 0.9000 ;
        RECT 0.1650 0.2550 0.4725 0.3300 ;
        RECT 0.3300 0.4050 0.4650 0.6450 ;
        RECT 0.0450 0.1500 0.1650 0.3300 ;
        RECT 0.5250 0.7200 0.6000 0.9000 ;
        RECT 0.4725 0.1575 0.5775 0.3300 ;
    END
END OR3_0011


MACRO OR3_0100
    CLASS CORE ;
    FOREIGN OR3_0100 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.7800 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 2.9925 0.2625 3.1500 0.3825 ;
        RECT 2.9925 0.6600 3.1500 0.7800 ;
        RECT 2.6775 0.2625 2.9925 0.7800 ;
        RECT 2.5200 0.2625 2.6775 0.3825 ;
        RECT 2.5200 0.6600 2.6775 0.7800 ;
        VIA 2.9925 0.3225 VIA12_slot ;
        VIA 2.9925 0.7200 VIA12_slot ;
        VIA 2.6775 0.3225 VIA12_slot ;
        VIA 2.6775 0.7200 VIA12_slot ;
        END
    END Z
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.4275 0.1125 0.8925 0.1875 ;
        RECT 0.4275 0.3975 0.4575 0.5475 ;
        RECT 0.3525 0.1125 0.4275 0.5475 ;
        VIA 0.4050 0.4725 VIA12_square ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.1925 0.5625 1.5075 0.6375 ;
        RECT 1.1175 0.4125 1.1925 0.6375 ;
        RECT 0.8025 0.4125 1.1175 0.4875 ;
        VIA 1.1550 0.4950 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.8225 0.5625 2.1375 0.6375 ;
        RECT 1.7475 0.4125 1.8225 0.6375 ;
        RECT 1.4325 0.4125 1.7475 0.4875 ;
        VIA 1.7850 0.4950 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 3.7125 -0.0750 3.7800 0.0750 ;
        RECT 3.6375 -0.0750 3.7125 0.2925 ;
        RECT 3.3150 -0.0750 3.6375 0.0750 ;
        RECT 3.1950 -0.0750 3.3150 0.1875 ;
        RECT 2.8950 -0.0750 3.1950 0.0750 ;
        RECT 2.7750 -0.0750 2.8950 0.1875 ;
        RECT 2.4750 -0.0750 2.7750 0.0750 ;
        RECT 2.3550 -0.0750 2.4750 0.1875 ;
        RECT 2.0550 -0.0750 2.3550 0.0750 ;
        RECT 1.9350 -0.0750 2.0550 0.1950 ;
        RECT 1.6350 -0.0750 1.9350 0.0750 ;
        RECT 1.5150 -0.0750 1.6350 0.1950 ;
        RECT 1.2150 -0.0750 1.5150 0.0750 ;
        RECT 1.0950 -0.0750 1.2150 0.1950 ;
        RECT 0.7950 -0.0750 1.0950 0.0750 ;
        RECT 0.6750 -0.0750 0.7950 0.1950 ;
        RECT 0.3750 -0.0750 0.6750 0.0750 ;
        RECT 0.2550 -0.0750 0.3750 0.1950 ;
        RECT 0.0000 -0.0750 0.2550 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 3.7125 0.9750 3.7800 1.1250 ;
        RECT 3.6375 0.6375 3.7125 1.1250 ;
        RECT 3.3150 0.9750 3.6375 1.1250 ;
        RECT 3.1950 0.8550 3.3150 1.1250 ;
        RECT 2.8950 0.9750 3.1950 1.1250 ;
        RECT 2.7750 0.8550 2.8950 1.1250 ;
        RECT 2.4750 0.9750 2.7750 1.1250 ;
        RECT 2.3550 0.8550 2.4750 1.1250 ;
        RECT 2.0325 0.9750 2.3550 1.1250 ;
        RECT 1.9575 0.6675 2.0325 1.1250 ;
        RECT 1.6350 0.9750 1.9575 1.1250 ;
        RECT 1.5150 0.7800 1.6350 1.1250 ;
        RECT 0.0000 0.9750 1.5150 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 3.6450 0.1875 3.7050 0.2475 ;
        RECT 3.6450 0.6675 3.7050 0.7275 ;
        RECT 3.6450 0.8325 3.7050 0.8925 ;
        RECT 3.5400 0.4650 3.6000 0.5250 ;
        RECT 3.4350 0.2850 3.4950 0.3450 ;
        RECT 3.4350 0.6900 3.4950 0.7500 ;
        RECT 3.3300 0.4650 3.3900 0.5250 ;
        RECT 3.2250 0.1275 3.2850 0.1875 ;
        RECT 3.2250 0.8625 3.2850 0.9225 ;
        RECT 3.1200 0.4650 3.1800 0.5250 ;
        RECT 3.0150 0.2850 3.0750 0.3450 ;
        RECT 3.0150 0.6900 3.0750 0.7500 ;
        RECT 2.9100 0.4650 2.9700 0.5250 ;
        RECT 2.8050 0.1275 2.8650 0.1875 ;
        RECT 2.8050 0.8625 2.8650 0.9225 ;
        RECT 2.7000 0.4650 2.7600 0.5250 ;
        RECT 2.5950 0.2850 2.6550 0.3450 ;
        RECT 2.5950 0.6900 2.6550 0.7500 ;
        RECT 2.4900 0.4650 2.5500 0.5250 ;
        RECT 2.3850 0.1275 2.4450 0.1875 ;
        RECT 2.3850 0.8625 2.4450 0.9225 ;
        RECT 2.2800 0.4650 2.3400 0.5250 ;
        RECT 2.1750 0.2925 2.2350 0.3525 ;
        RECT 2.1750 0.6900 2.2350 0.7500 ;
        RECT 2.0700 0.4650 2.1300 0.5250 ;
        RECT 1.9650 0.1275 2.0250 0.1875 ;
        RECT 1.9650 0.6975 2.0250 0.7575 ;
        RECT 1.9650 0.8625 2.0250 0.9225 ;
        RECT 1.8600 0.4650 1.9200 0.5250 ;
        RECT 1.7550 0.1725 1.8150 0.2325 ;
        RECT 1.7550 0.6450 1.8150 0.7050 ;
        RECT 1.7550 0.8325 1.8150 0.8925 ;
        RECT 1.6500 0.4650 1.7100 0.5250 ;
        RECT 1.5450 0.1275 1.6050 0.1875 ;
        RECT 1.5450 0.8025 1.6050 0.8625 ;
        RECT 1.4400 0.4650 1.5000 0.5250 ;
        RECT 1.3350 0.1725 1.3950 0.2325 ;
        RECT 1.3350 0.6450 1.3950 0.7050 ;
        RECT 1.3350 0.8325 1.3950 0.8925 ;
        RECT 1.2300 0.4650 1.2900 0.5250 ;
        RECT 1.1250 0.1275 1.1850 0.1875 ;
        RECT 1.1250 0.8025 1.1850 0.8625 ;
        RECT 1.0200 0.4650 1.0800 0.5250 ;
        RECT 0.9150 0.1725 0.9750 0.2325 ;
        RECT 0.9150 0.6675 0.9750 0.7275 ;
        RECT 0.8100 0.4650 0.8700 0.5250 ;
        RECT 0.7050 0.1275 0.7650 0.1875 ;
        RECT 0.7050 0.6675 0.7650 0.7275 ;
        RECT 0.7050 0.8325 0.7650 0.8925 ;
        RECT 0.6000 0.4650 0.6600 0.5250 ;
        RECT 0.4950 0.2775 0.5550 0.3375 ;
        RECT 0.4950 0.6525 0.5550 0.7125 ;
        RECT 0.3900 0.4650 0.4500 0.5250 ;
        RECT 0.2850 0.1275 0.3450 0.1875 ;
        RECT 0.2850 0.8025 0.3450 0.8625 ;
        RECT 0.1800 0.4650 0.2400 0.5250 ;
        RECT 0.0750 0.2625 0.1350 0.3225 ;
        RECT 0.0750 0.6525 0.1350 0.7125 ;
        RECT 0.0750 0.8175 0.1350 0.8775 ;
        LAYER M1 ;
        RECT 2.1000 0.4575 3.6300 0.5325 ;
        RECT 2.1750 0.2625 3.5175 0.3825 ;
        RECT 2.1525 0.6600 3.5175 0.7800 ;
        RECT 2.0250 0.2700 2.1000 0.5325 ;
        RECT 1.8375 0.2700 2.0250 0.3450 ;
        RECT 1.4100 0.4350 1.9500 0.5400 ;
        RECT 1.7250 0.6150 1.8450 0.9000 ;
        RECT 1.7325 0.1500 1.8375 0.3450 ;
        RECT 1.4175 0.2700 1.7325 0.3450 ;
        RECT 1.4250 0.6150 1.7250 0.6975 ;
        RECT 1.3050 0.6150 1.4250 0.8925 ;
        RECT 1.3125 0.1500 1.4175 0.3450 ;
        RECT 0.7800 0.4350 1.3200 0.5400 ;
        RECT 0.9975 0.2700 1.3125 0.3450 ;
        RECT 0.9975 0.6150 1.3050 0.6975 ;
        RECT 1.0950 0.7725 1.2150 0.9000 ;
        RECT 0.7875 0.8250 1.0950 0.9000 ;
        RECT 0.8925 0.1500 0.9975 0.3450 ;
        RECT 0.8925 0.6150 0.9975 0.7500 ;
        RECT 0.1575 0.2700 0.8925 0.3450 ;
        RECT 0.6825 0.6450 0.7875 0.9000 ;
        RECT 0.1500 0.4350 0.6900 0.5400 ;
        RECT 0.3750 0.8250 0.6825 0.9000 ;
        RECT 0.4575 0.6150 0.6075 0.7275 ;
        RECT 0.1575 0.6150 0.4575 0.6900 ;
        RECT 0.2550 0.7725 0.3750 0.9000 ;
        RECT 0.0525 0.2400 0.1575 0.3450 ;
        RECT 0.0525 0.6150 0.1575 0.9000 ;
        LAYER VIA1 ;
        RECT 0.5925 0.2700 0.6675 0.3450 ;
        RECT 0.4950 0.6300 0.5700 0.7050 ;
        LAYER M2 ;
        RECT 3.0225 0.2625 3.1500 0.3825 ;
        RECT 3.0225 0.6600 3.1500 0.7800 ;
        RECT 2.5200 0.2625 2.6475 0.3825 ;
        RECT 2.5200 0.6600 2.6475 0.7800 ;
        RECT 0.6225 0.2700 0.7425 0.3450 ;
        RECT 0.5475 0.2700 0.6225 0.7050 ;
        RECT 0.4500 0.6300 0.5475 0.7050 ;
    END
END OR3_0100


MACRO OR3_0111
    CLASS CORE ;
    FOREIGN OR3_0111 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.3100 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 1.6275 0.2625 1.9425 0.7275 ;
        VIA 1.7850 0.3225 VIA12_slot ;
        VIA 1.7850 0.6675 VIA12_slot ;
        END
    END Z
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.7875 0.4125 1.0125 0.4875 ;
        RECT 0.6825 0.4125 0.7875 0.5625 ;
        RECT 0.5475 0.4125 0.6825 0.4875 ;
        VIA 0.7350 0.4875 VIA12_square ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.9975 0.7125 1.4625 0.7875 ;
        RECT 0.8925 0.6000 0.9975 0.7875 ;
        VIA 0.9450 0.6750 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.2300 0.4200 1.2600 0.5850 ;
        RECT 1.1550 0.2625 1.2300 0.5850 ;
        RECT 0.4275 0.2625 1.1550 0.3375 ;
        RECT 0.3525 0.2625 0.4275 0.6375 ;
        RECT 0.1650 0.5625 0.3525 0.6375 ;
        VIA 1.2075 0.5025 VIA12_square ;
        VIA 0.2775 0.6000 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 2.2425 -0.0750 2.3100 0.0750 ;
        RECT 2.1675 -0.0750 2.2425 0.3150 ;
        RECT 1.8450 -0.0750 2.1675 0.0750 ;
        RECT 1.7250 -0.0750 1.8450 0.1950 ;
        RECT 1.4250 -0.0750 1.7250 0.0750 ;
        RECT 1.3050 -0.0750 1.4250 0.1950 ;
        RECT 1.0050 -0.0750 1.3050 0.0750 ;
        RECT 0.8850 -0.0750 1.0050 0.1950 ;
        RECT 0.5850 -0.0750 0.8850 0.0750 ;
        RECT 0.4650 -0.0750 0.5850 0.1950 ;
        RECT 0.1425 -0.0750 0.4650 0.0750 ;
        RECT 0.0675 -0.0750 0.1425 0.2625 ;
        RECT 0.0000 -0.0750 0.0675 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 2.2425 0.9750 2.3100 1.1250 ;
        RECT 2.1675 0.6375 2.2425 1.1250 ;
        RECT 1.8225 0.9750 2.1675 1.1250 ;
        RECT 1.7475 0.8175 1.8225 1.1250 ;
        RECT 1.4250 0.9750 1.7475 1.1250 ;
        RECT 1.3050 0.8550 1.4250 1.1250 ;
        RECT 0.1575 0.9750 1.3050 1.1250 ;
        RECT 0.0525 0.6450 0.1575 1.1250 ;
        RECT 0.0000 0.9750 0.0525 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 2.1750 0.2250 2.2350 0.2850 ;
        RECT 2.1750 0.6675 2.2350 0.7275 ;
        RECT 2.1750 0.8325 2.2350 0.8925 ;
        RECT 2.0700 0.4650 2.1300 0.5250 ;
        RECT 1.9650 0.2250 2.0250 0.2850 ;
        RECT 1.9650 0.7575 2.0250 0.8175 ;
        RECT 1.8600 0.4650 1.9200 0.5250 ;
        RECT 1.7550 0.1275 1.8150 0.1875 ;
        RECT 1.7550 0.8475 1.8150 0.9075 ;
        RECT 1.6500 0.4650 1.7100 0.5250 ;
        RECT 1.5450 0.2250 1.6050 0.2850 ;
        RECT 1.5450 0.7575 1.6050 0.8175 ;
        RECT 1.4400 0.4650 1.5000 0.5250 ;
        RECT 1.3350 0.1275 1.3950 0.1875 ;
        RECT 1.3350 0.8625 1.3950 0.9225 ;
        RECT 1.2300 0.4800 1.2900 0.5400 ;
        RECT 1.1250 0.1725 1.1850 0.2325 ;
        RECT 1.0200 0.4800 1.0800 0.5400 ;
        RECT 0.9150 0.1275 0.9750 0.1875 ;
        RECT 0.8100 0.4650 0.8700 0.5250 ;
        RECT 0.7050 0.1725 0.7650 0.2325 ;
        RECT 0.7050 0.8175 0.7650 0.8775 ;
        RECT 0.6000 0.4650 0.6600 0.5250 ;
        RECT 0.4950 0.1275 0.5550 0.1875 ;
        RECT 0.3900 0.4875 0.4500 0.5475 ;
        RECT 0.2850 0.1725 0.3450 0.2325 ;
        RECT 0.1800 0.4725 0.2400 0.5325 ;
        RECT 0.0750 0.1575 0.1350 0.2175 ;
        RECT 0.0750 0.6675 0.1350 0.7275 ;
        RECT 0.0750 0.8325 0.1350 0.8925 ;
        LAYER M1 ;
        RECT 1.4625 0.4425 2.1600 0.5475 ;
        RECT 1.9425 0.1950 2.0475 0.3675 ;
        RECT 1.9575 0.6225 2.0325 0.8700 ;
        RECT 1.6125 0.6225 1.9575 0.7125 ;
        RECT 1.6275 0.2775 1.9425 0.3675 ;
        RECT 1.5375 0.1950 1.6275 0.3675 ;
        RECT 1.5375 0.6225 1.6125 0.8700 ;
        RECT 1.3875 0.2700 1.4625 0.7800 ;
        RECT 1.2075 0.2700 1.3875 0.3450 ;
        RECT 1.2300 0.7050 1.3875 0.7800 ;
        RECT 1.1550 0.4200 1.3050 0.6300 ;
        RECT 1.1550 0.7050 1.2300 0.8850 ;
        RECT 1.1025 0.1500 1.2075 0.3450 ;
        RECT 0.6675 0.8100 1.1550 0.8850 ;
        RECT 0.7875 0.2700 1.1025 0.3450 ;
        RECT 1.0050 0.4500 1.0800 0.7125 ;
        RECT 0.4650 0.6375 1.0050 0.7125 ;
        RECT 0.5925 0.4350 0.8775 0.5625 ;
        RECT 0.6825 0.1500 0.7875 0.3450 ;
        RECT 0.3675 0.2700 0.6825 0.3450 ;
        RECT 0.3900 0.4500 0.4650 0.7125 ;
        RECT 0.2625 0.1500 0.3675 0.3450 ;
        RECT 0.2400 0.4200 0.3150 0.7125 ;
        RECT 0.1050 0.4200 0.2400 0.5550 ;
    END
END OR3_0111


MACRO OR3_1000
    CLASS CORE ;
    FOREIGN OR3_1000 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.0500 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.9375 0.1500 1.0125 0.9000 ;
        RECT 0.8850 0.1500 0.9375 0.3825 ;
        RECT 0.8925 0.6675 0.9375 0.9000 ;
        END
    END Z
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.1350 0.5625 0.6000 0.6375 ;
        VIA 0.2475 0.6000 VIA12_square ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.4500 0.8625 0.9150 0.9375 ;
        RECT 0.3450 0.7650 0.4500 0.9375 ;
        VIA 0.3975 0.8475 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.3525 0.4125 0.8175 0.4875 ;
        VIA 0.5775 0.4500 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.7950 -0.0750 1.0500 0.0750 ;
        RECT 0.6750 -0.0750 0.7950 0.1800 ;
        RECT 0.3750 -0.0750 0.6750 0.0750 ;
        RECT 0.2550 -0.0750 0.3750 0.1800 ;
        RECT 0.0000 -0.0750 0.2550 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.7950 0.9750 1.0500 1.1250 ;
        RECT 0.6750 0.8700 0.7950 1.1250 ;
        RECT 0.0000 0.9750 0.6750 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 0.9150 0.1575 0.9750 0.2175 ;
        RECT 0.9150 0.8175 0.9750 0.8775 ;
        RECT 0.8025 0.4950 0.8625 0.5550 ;
        RECT 0.7050 0.1200 0.7650 0.1800 ;
        RECT 0.7050 0.8700 0.7650 0.9300 ;
        RECT 0.6000 0.4875 0.6600 0.5475 ;
        RECT 0.4950 0.1725 0.5550 0.2325 ;
        RECT 0.3825 0.6375 0.4425 0.6975 ;
        RECT 0.2850 0.1200 0.3450 0.1800 ;
        RECT 0.1875 0.4950 0.2475 0.5550 ;
        RECT 0.0750 0.1575 0.1350 0.2175 ;
        RECT 0.0750 0.8175 0.1350 0.8775 ;
        LAYER M1 ;
        RECT 0.8100 0.4650 0.8625 0.5850 ;
        RECT 0.7350 0.2550 0.8100 0.5850 ;
        RECT 0.5775 0.2550 0.7350 0.3300 ;
        RECT 0.5175 0.4050 0.6600 0.6450 ;
        RECT 0.4725 0.1500 0.5775 0.3300 ;
        RECT 0.4950 0.4050 0.5175 0.5100 ;
        RECT 0.4425 0.8025 0.5100 0.8925 ;
        RECT 0.1650 0.2550 0.4725 0.3300 ;
        RECT 0.3675 0.6075 0.4425 0.8925 ;
        RECT 0.2850 0.8025 0.3675 0.8925 ;
        RECT 0.1875 0.4050 0.2925 0.7050 ;
        RECT 0.1125 0.1500 0.1650 0.3300 ;
        RECT 0.1125 0.7950 0.1575 0.9000 ;
        RECT 0.0375 0.1500 0.1125 0.9000 ;
    END
END OR3_1000


MACRO OR3_1010
    CLASS CORE ;
    FOREIGN OR3_1010 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.0500 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.9375 0.2175 1.0125 0.8325 ;
        RECT 0.9150 0.2175 0.9375 0.3825 ;
        RECT 0.9075 0.6675 0.9375 0.8325 ;
        END
    END Z
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.1350 0.5625 0.6000 0.6375 ;
        VIA 0.2475 0.6000 VIA12_square ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.4500 0.8625 0.9150 0.9375 ;
        RECT 0.3450 0.7650 0.4500 0.9375 ;
        VIA 0.3975 0.8475 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.3525 0.4125 0.8175 0.4875 ;
        VIA 0.6000 0.4500 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.7950 -0.0750 1.0500 0.0750 ;
        RECT 0.6750 -0.0750 0.7950 0.1800 ;
        RECT 0.3750 -0.0750 0.6750 0.0750 ;
        RECT 0.2550 -0.0750 0.3750 0.1800 ;
        RECT 0.0000 -0.0750 0.2550 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.7950 0.9750 1.0500 1.1250 ;
        RECT 0.6750 0.8700 0.7950 1.1250 ;
        RECT 0.0000 0.9750 0.6750 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 0.9150 0.2775 0.9750 0.3375 ;
        RECT 0.9150 0.7425 0.9750 0.8025 ;
        RECT 0.8025 0.4950 0.8625 0.5550 ;
        RECT 0.7050 0.1200 0.7650 0.1800 ;
        RECT 0.7050 0.8700 0.7650 0.9300 ;
        RECT 0.6000 0.4875 0.6600 0.5475 ;
        RECT 0.4950 0.1725 0.5550 0.2325 ;
        RECT 0.3825 0.4875 0.4425 0.5475 ;
        RECT 0.2850 0.1200 0.3450 0.1800 ;
        RECT 0.1875 0.4950 0.2475 0.5550 ;
        RECT 0.0750 0.1725 0.1350 0.2325 ;
        RECT 0.0750 0.7950 0.1350 0.8550 ;
        LAYER M1 ;
        RECT 0.8325 0.4650 0.8625 0.5850 ;
        RECT 0.7575 0.2550 0.8325 0.5850 ;
        RECT 0.5775 0.2550 0.7575 0.3300 ;
        RECT 0.5175 0.4050 0.6825 0.6450 ;
        RECT 0.4725 0.1500 0.5775 0.3300 ;
        RECT 0.4425 0.8025 0.5100 0.8925 ;
        RECT 0.1575 0.2550 0.4725 0.3300 ;
        RECT 0.3675 0.4350 0.4425 0.8925 ;
        RECT 0.2850 0.8025 0.3675 0.8925 ;
        RECT 0.1875 0.4050 0.2925 0.7050 ;
        RECT 0.1125 0.1500 0.1575 0.3300 ;
        RECT 0.1125 0.7650 0.1425 0.8850 ;
        RECT 0.0375 0.1500 0.1125 0.8850 ;
    END
END OR3_1010


MACRO OR4_0011
    CLASS CORE ;
    FOREIGN OR4_0011 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.4700 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 1.3575 0.3075 1.4325 0.7350 ;
        RECT 1.1925 0.3075 1.3575 0.3825 ;
        RECT 1.1925 0.6600 1.3575 0.7350 ;
        RECT 1.1175 0.2175 1.1925 0.3825 ;
        RECT 1.1175 0.6600 1.1925 0.8325 ;
        END
    END Z
    PIN A4
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1425 0.4500 0.2400 0.6375 ;
        RECT 0.0675 0.3675 0.1425 0.6375 ;
        END
    END A4
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.4575 0.8625 0.9225 0.9375 ;
        RECT 0.4575 0.4875 0.4875 0.6450 ;
        RECT 0.3825 0.4875 0.4575 0.9375 ;
        VIA 0.4350 0.5625 VIA12_square ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.6825 0.7125 1.1175 0.7875 ;
        RECT 0.5775 0.4800 0.6825 0.7875 ;
        VIA 0.6300 0.5625 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.8925 0.4650 0.9225 0.5700 ;
        RECT 0.8175 0.2625 0.8925 0.5700 ;
        RECT 0.3525 0.2625 0.8175 0.3375 ;
        VIA 0.8550 0.4875 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.4250 -0.0750 1.4700 0.0750 ;
        RECT 1.3050 -0.0750 1.4250 0.2325 ;
        RECT 1.0050 -0.0750 1.3050 0.0750 ;
        RECT 0.8850 -0.0750 1.0050 0.1800 ;
        RECT 0.5850 -0.0750 0.8850 0.0750 ;
        RECT 0.4650 -0.0750 0.5850 0.1800 ;
        RECT 0.1425 -0.0750 0.4650 0.0750 ;
        RECT 0.0675 -0.0750 0.1425 0.2625 ;
        RECT 0.0000 -0.0750 0.0675 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.4175 0.9750 1.4700 1.1250 ;
        RECT 1.3125 0.8100 1.4175 1.1250 ;
        RECT 1.0050 0.9750 1.3125 1.1250 ;
        RECT 0.8850 0.8700 1.0050 1.1250 ;
        RECT 0.0000 0.9750 0.8850 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.3350 0.1650 1.3950 0.2250 ;
        RECT 1.3350 0.8325 1.3950 0.8925 ;
        RECT 1.2225 0.4875 1.2825 0.5475 ;
        RECT 1.1250 0.2700 1.1850 0.3300 ;
        RECT 1.1250 0.7200 1.1850 0.7800 ;
        RECT 1.0200 0.4875 1.0800 0.5475 ;
        RECT 0.9150 0.1200 0.9750 0.1800 ;
        RECT 0.9150 0.8700 0.9750 0.9300 ;
        RECT 0.8100 0.4725 0.8700 0.5325 ;
        RECT 0.7050 0.2625 0.7650 0.3225 ;
        RECT 0.6000 0.4800 0.6600 0.5400 ;
        RECT 0.4950 0.1200 0.5550 0.1800 ;
        RECT 0.3900 0.4800 0.4500 0.5400 ;
        RECT 0.2850 0.1950 0.3450 0.2550 ;
        RECT 0.1800 0.4950 0.2400 0.5550 ;
        RECT 0.0750 0.1650 0.1350 0.2250 ;
        RECT 0.0750 0.7875 0.1350 0.8475 ;
        LAYER M1 ;
        RECT 1.0425 0.4575 1.2825 0.5775 ;
        RECT 0.9675 0.2550 1.0425 0.7950 ;
        RECT 0.3675 0.2550 0.9675 0.3300 ;
        RECT 0.1425 0.7200 0.9675 0.7950 ;
        RECT 0.7575 0.4050 0.8925 0.6450 ;
        RECT 0.5475 0.4050 0.6825 0.6450 ;
        RECT 0.3300 0.4050 0.4725 0.6450 ;
        RECT 0.2625 0.1650 0.3675 0.3300 ;
        RECT 0.0675 0.7200 0.1425 0.8850 ;
    END
END OR4_0011


MACRO OR4_0100
    CLASS CORE ;
    FOREIGN OR4_0100 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.4100 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 3.6225 0.2625 3.7800 0.3825 ;
        RECT 3.6225 0.6600 3.7800 0.7800 ;
        RECT 3.3075 0.2625 3.6225 0.7800 ;
        RECT 3.1500 0.2625 3.3075 0.3825 ;
        RECT 3.1500 0.6600 3.3075 0.7800 ;
        VIA 3.6225 0.3225 VIA12_slot ;
        VIA 3.6225 0.7200 VIA12_slot ;
        VIA 3.3075 0.3225 VIA12_slot ;
        VIA 3.3075 0.7200 VIA12_slot ;
        END
    END Z
    PIN A4
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.5025 0.1125 0.9675 0.1875 ;
        RECT 0.4275 0.1125 0.5025 0.5700 ;
        RECT 0.3525 0.4650 0.4275 0.5700 ;
        VIA 0.4275 0.5175 VIA12_square ;
        END
    END A4
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.1925 0.5625 1.5075 0.6375 ;
        RECT 1.1175 0.4125 1.1925 0.6375 ;
        RECT 0.8025 0.4125 1.1175 0.4875 ;
        VIA 1.1550 0.5175 VIA12_square ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.8225 0.5625 2.1375 0.6375 ;
        RECT 1.7475 0.4125 1.8225 0.6375 ;
        RECT 1.4325 0.4125 1.7475 0.4875 ;
        VIA 1.7850 0.5175 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 2.4525 0.5625 2.7675 0.6375 ;
        RECT 2.3775 0.4125 2.4525 0.6375 ;
        RECT 2.0625 0.4125 2.3775 0.4875 ;
        VIA 2.4150 0.5325 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 4.3425 -0.0750 4.4100 0.0750 ;
        RECT 4.2675 -0.0750 4.3425 0.2925 ;
        RECT 3.9450 -0.0750 4.2675 0.0750 ;
        RECT 3.8250 -0.0750 3.9450 0.1875 ;
        RECT 3.5250 -0.0750 3.8250 0.0750 ;
        RECT 3.4050 -0.0750 3.5250 0.1875 ;
        RECT 3.1050 -0.0750 3.4050 0.0750 ;
        RECT 2.9850 -0.0750 3.1050 0.1875 ;
        RECT 2.6850 -0.0750 2.9850 0.0750 ;
        RECT 2.5650 -0.0750 2.6850 0.2325 ;
        RECT 2.2650 -0.0750 2.5650 0.0750 ;
        RECT 2.1450 -0.0750 2.2650 0.2325 ;
        RECT 1.8450 -0.0750 2.1450 0.0750 ;
        RECT 1.7250 -0.0750 1.8450 0.2325 ;
        RECT 1.4250 -0.0750 1.7250 0.0750 ;
        RECT 1.3050 -0.0750 1.4250 0.2325 ;
        RECT 1.0050 -0.0750 1.3050 0.0750 ;
        RECT 0.8850 -0.0750 1.0050 0.2325 ;
        RECT 0.5850 -0.0750 0.8850 0.0750 ;
        RECT 0.4650 -0.0750 0.5850 0.2325 ;
        RECT 0.1425 -0.0750 0.4650 0.0750 ;
        RECT 0.0675 -0.0750 0.1425 0.2475 ;
        RECT 0.0000 -0.0750 0.0675 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 4.3575 0.9750 4.4100 1.1250 ;
        RECT 4.2525 0.6450 4.3575 1.1250 ;
        RECT 3.9450 0.9750 4.2525 1.1250 ;
        RECT 3.8250 0.8550 3.9450 1.1250 ;
        RECT 3.5250 0.9750 3.8250 1.1250 ;
        RECT 3.4050 0.8550 3.5250 1.1250 ;
        RECT 3.1050 0.9750 3.4050 1.1250 ;
        RECT 2.9850 0.8550 3.1050 1.1250 ;
        RECT 2.6850 0.9750 2.9850 1.1250 ;
        RECT 2.5800 0.6750 2.6850 1.1250 ;
        RECT 2.2575 0.9750 2.5800 1.1250 ;
        RECT 2.1525 0.8250 2.2575 1.1250 ;
        RECT 0.0000 0.9750 2.1525 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 4.2750 0.1875 4.3350 0.2475 ;
        RECT 4.2750 0.6675 4.3350 0.7275 ;
        RECT 4.2750 0.8325 4.3350 0.8925 ;
        RECT 4.1700 0.4800 4.2300 0.5400 ;
        RECT 4.0650 0.2850 4.1250 0.3450 ;
        RECT 4.0650 0.6900 4.1250 0.7500 ;
        RECT 3.9600 0.4800 4.0200 0.5400 ;
        RECT 3.8550 0.1275 3.9150 0.1875 ;
        RECT 3.8550 0.8625 3.9150 0.9225 ;
        RECT 3.7500 0.4800 3.8100 0.5400 ;
        RECT 3.6450 0.2850 3.7050 0.3450 ;
        RECT 3.6450 0.6900 3.7050 0.7500 ;
        RECT 3.5400 0.4800 3.6000 0.5400 ;
        RECT 3.4350 0.1275 3.4950 0.1875 ;
        RECT 3.4350 0.8625 3.4950 0.9225 ;
        RECT 3.3300 0.4800 3.3900 0.5400 ;
        RECT 3.2250 0.2850 3.2850 0.3450 ;
        RECT 3.2250 0.6900 3.2850 0.7500 ;
        RECT 3.1200 0.4800 3.1800 0.5400 ;
        RECT 3.0150 0.1275 3.0750 0.1875 ;
        RECT 3.0150 0.8625 3.0750 0.9225 ;
        RECT 2.9100 0.4800 2.9700 0.5400 ;
        RECT 2.8050 0.2850 2.8650 0.3450 ;
        RECT 2.8050 0.6900 2.8650 0.7500 ;
        RECT 2.7000 0.4800 2.7600 0.5400 ;
        RECT 2.5950 0.1575 2.6550 0.2175 ;
        RECT 2.5950 0.7050 2.6550 0.7650 ;
        RECT 2.5950 0.8700 2.6550 0.9300 ;
        RECT 2.4900 0.4950 2.5500 0.5550 ;
        RECT 2.3850 0.3150 2.4450 0.3750 ;
        RECT 2.3850 0.6825 2.4450 0.7425 ;
        RECT 2.2800 0.4950 2.3400 0.5550 ;
        RECT 2.1750 0.1575 2.2350 0.2175 ;
        RECT 2.1750 0.8475 2.2350 0.9075 ;
        RECT 2.0700 0.4950 2.1300 0.5550 ;
        RECT 1.9650 0.3150 2.0250 0.3750 ;
        RECT 1.9650 0.6825 2.0250 0.7425 ;
        RECT 1.8600 0.4875 1.9200 0.5475 ;
        RECT 1.7550 0.1575 1.8150 0.2175 ;
        RECT 1.7550 0.8325 1.8150 0.8925 ;
        RECT 1.6500 0.4875 1.7100 0.5475 ;
        RECT 1.5450 0.3150 1.6050 0.3750 ;
        RECT 1.5450 0.6825 1.6050 0.7425 ;
        RECT 1.4400 0.4875 1.5000 0.5475 ;
        RECT 1.3350 0.1575 1.3950 0.2175 ;
        RECT 1.3350 0.8325 1.3950 0.8925 ;
        RECT 1.2300 0.4875 1.2900 0.5475 ;
        RECT 1.1250 0.3150 1.1850 0.3750 ;
        RECT 1.1250 0.6825 1.1850 0.7425 ;
        RECT 1.0200 0.4875 1.0800 0.5475 ;
        RECT 0.9150 0.1575 0.9750 0.2175 ;
        RECT 0.9150 0.8325 0.9750 0.8925 ;
        RECT 0.8100 0.4875 0.8700 0.5475 ;
        RECT 0.7050 0.3150 0.7650 0.3750 ;
        RECT 0.7050 0.7575 0.7650 0.8175 ;
        RECT 0.6000 0.4875 0.6600 0.5475 ;
        RECT 0.4950 0.1575 0.5550 0.2175 ;
        RECT 0.4950 0.6825 0.5550 0.7425 ;
        RECT 0.3900 0.4875 0.4500 0.5475 ;
        RECT 0.2850 0.2775 0.3450 0.3375 ;
        RECT 0.2850 0.8325 0.3450 0.8925 ;
        RECT 0.1800 0.4875 0.2400 0.5475 ;
        RECT 0.0750 0.1575 0.1350 0.2175 ;
        RECT 0.0750 0.6975 0.1350 0.7575 ;
        LAYER M1 ;
        RECT 2.7075 0.4725 4.2600 0.5475 ;
        RECT 2.7825 0.2625 4.1475 0.3825 ;
        RECT 2.7825 0.6600 4.1475 0.7800 ;
        RECT 2.6325 0.3075 2.7075 0.5475 ;
        RECT 0.3675 0.3075 2.6325 0.3900 ;
        RECT 2.0325 0.4650 2.5575 0.5850 ;
        RECT 1.5150 0.6750 2.4750 0.7500 ;
        RECT 1.4025 0.4650 1.9575 0.5700 ;
        RECT 0.8850 0.8250 1.8450 0.9000 ;
        RECT 0.7725 0.4650 1.3275 0.5700 ;
        RECT 0.7725 0.6750 1.2150 0.7500 ;
        RECT 0.6975 0.6750 0.7725 0.9000 ;
        RECT 0.1500 0.4650 0.6975 0.5700 ;
        RECT 0.2550 0.8250 0.6975 0.9000 ;
        RECT 0.1575 0.6750 0.5925 0.7500 ;
        RECT 0.2625 0.2400 0.3675 0.3900 ;
        RECT 0.0525 0.6750 0.1575 0.7800 ;
        LAYER VIA1 ;
        RECT 0.5925 0.3150 0.6675 0.3900 ;
        RECT 0.4725 0.6750 0.5475 0.7500 ;
        LAYER M2 ;
        RECT 3.6525 0.2625 3.7800 0.3825 ;
        RECT 3.6525 0.6600 3.7800 0.7800 ;
        RECT 3.1500 0.2625 3.2775 0.3825 ;
        RECT 3.1500 0.6600 3.2775 0.7800 ;
        RECT 0.5775 0.2775 0.6825 0.7650 ;
        RECT 0.4350 0.6600 0.5775 0.7650 ;
    END
END OR4_0100


MACRO OR4_0111
    CLASS CORE ;
    FOREIGN OR4_0111 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.7300 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 2.0475 0.2625 2.3625 0.7275 ;
        VIA 2.2050 0.3225 VIA12_slot ;
        VIA 2.2050 0.6675 VIA12_slot ;
        END
    END Z
    PIN A4
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.0200 0.4125 1.2375 0.4875 ;
        RECT 0.8700 0.4125 1.0200 0.5625 ;
        RECT 0.6975 0.4125 0.8700 0.4875 ;
        VIA 0.9450 0.5100 VIA12_square ;
        END
    END A4
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.7875 0.7125 1.2525 0.7875 ;
        RECT 0.6825 0.6375 0.7875 0.7875 ;
        VIA 0.7350 0.7125 VIA12_square ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.4325 0.4800 1.4625 0.6450 ;
        RECT 1.3575 0.2625 1.4325 0.6450 ;
        RECT 0.5775 0.2625 1.3575 0.3375 ;
        RECT 0.5025 0.2625 0.5775 0.7875 ;
        RECT 0.3675 0.7125 0.5025 0.7875 ;
        VIA 1.4100 0.5625 VIA12_square ;
        VIA 0.4800 0.7500 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.6425 0.4800 1.6725 0.6450 ;
        RECT 1.5675 0.1125 1.6425 0.6450 ;
        RECT 0.4275 0.1125 1.5675 0.1875 ;
        RECT 0.3525 0.1125 0.4275 0.6375 ;
        RECT 0.1575 0.5625 0.3525 0.6375 ;
        VIA 1.6200 0.5625 VIA12_square ;
        VIA 0.2700 0.6000 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 2.6625 -0.0750 2.7300 0.0750 ;
        RECT 2.5875 -0.0750 2.6625 0.3150 ;
        RECT 2.2650 -0.0750 2.5875 0.0750 ;
        RECT 2.1450 -0.0750 2.2650 0.1950 ;
        RECT 1.8450 -0.0750 2.1450 0.0750 ;
        RECT 1.7250 -0.0750 1.8450 0.2325 ;
        RECT 1.4250 -0.0750 1.7250 0.0750 ;
        RECT 1.3050 -0.0750 1.4250 0.2325 ;
        RECT 1.0050 -0.0750 1.3050 0.0750 ;
        RECT 0.8850 -0.0750 1.0050 0.2325 ;
        RECT 0.5850 -0.0750 0.8850 0.0750 ;
        RECT 0.4650 -0.0750 0.5850 0.2325 ;
        RECT 0.1500 -0.0750 0.4650 0.0750 ;
        RECT 0.0600 -0.0750 0.1500 0.3075 ;
        RECT 0.0000 -0.0750 0.0600 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 2.6775 0.9750 2.7300 1.1250 ;
        RECT 2.5725 0.6450 2.6775 1.1250 ;
        RECT 2.2425 0.9750 2.5725 1.1250 ;
        RECT 2.1675 0.8175 2.2425 1.1250 ;
        RECT 1.8375 0.9750 2.1675 1.1250 ;
        RECT 1.7325 0.8025 1.8375 1.1250 ;
        RECT 0.1575 0.9750 1.7325 1.1250 ;
        RECT 0.0525 0.6450 0.1575 1.1250 ;
        RECT 0.0000 0.9750 0.0525 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 2.5950 0.2250 2.6550 0.2850 ;
        RECT 2.5950 0.6675 2.6550 0.7275 ;
        RECT 2.5950 0.8325 2.6550 0.8925 ;
        RECT 2.4900 0.4650 2.5500 0.5250 ;
        RECT 2.3850 0.2250 2.4450 0.2850 ;
        RECT 2.3850 0.7575 2.4450 0.8175 ;
        RECT 2.2800 0.4650 2.3400 0.5250 ;
        RECT 2.1750 0.1275 2.2350 0.1875 ;
        RECT 2.1750 0.8475 2.2350 0.9075 ;
        RECT 2.0700 0.4650 2.1300 0.5250 ;
        RECT 1.9650 0.2250 2.0250 0.2850 ;
        RECT 1.9650 0.7575 2.0250 0.8175 ;
        RECT 1.8600 0.4650 1.9200 0.5250 ;
        RECT 1.7550 0.1575 1.8150 0.2175 ;
        RECT 1.7550 0.8250 1.8150 0.8850 ;
        RECT 1.6500 0.4950 1.7100 0.5550 ;
        RECT 1.5450 0.3150 1.6050 0.3750 ;
        RECT 1.4400 0.4950 1.5000 0.5550 ;
        RECT 1.3350 0.1575 1.3950 0.2175 ;
        RECT 1.2300 0.4950 1.2900 0.5550 ;
        RECT 1.1250 0.3150 1.1850 0.3750 ;
        RECT 1.0200 0.4950 1.0800 0.5550 ;
        RECT 0.9150 0.1575 0.9750 0.2175 ;
        RECT 0.9150 0.8325 0.9750 0.8925 ;
        RECT 0.8100 0.4950 0.8700 0.5550 ;
        RECT 0.7050 0.3150 0.7650 0.3750 ;
        RECT 0.6000 0.4950 0.6600 0.5550 ;
        RECT 0.4950 0.1575 0.5550 0.2175 ;
        RECT 0.3900 0.4950 0.4500 0.5550 ;
        RECT 0.2850 0.2775 0.3450 0.3375 ;
        RECT 0.1800 0.4875 0.2400 0.5475 ;
        RECT 0.0750 0.2100 0.1350 0.2700 ;
        RECT 0.0750 0.6675 0.1350 0.7275 ;
        RECT 0.0750 0.8325 0.1350 0.8925 ;
        LAYER M1 ;
        RECT 1.8675 0.4500 2.5800 0.5400 ;
        RECT 2.3625 0.1950 2.4675 0.3675 ;
        RECT 2.3775 0.6225 2.4525 0.8700 ;
        RECT 2.0325 0.6225 2.3775 0.7125 ;
        RECT 2.0475 0.2775 2.3625 0.3675 ;
        RECT 1.9425 0.1950 2.0475 0.3675 ;
        RECT 1.9575 0.6225 2.0325 0.8700 ;
        RECT 1.7925 0.3075 1.8675 0.5400 ;
        RECT 0.3675 0.3075 1.7925 0.3900 ;
        RECT 1.5825 0.4650 1.7175 0.7050 ;
        RECT 1.4925 0.7950 1.6575 0.9000 ;
        RECT 1.3725 0.4650 1.5075 0.7050 ;
        RECT 0.8850 0.8250 1.4925 0.9000 ;
        RECT 1.1925 0.4650 1.2975 0.7500 ;
        RECT 0.7125 0.6750 1.1925 0.7500 ;
        RECT 0.8025 0.4650 1.0875 0.6000 ;
        RECT 0.6375 0.4725 0.7125 0.7500 ;
        RECT 0.5775 0.4725 0.6375 0.5775 ;
        RECT 0.5025 0.6600 0.5625 0.8250 ;
        RECT 0.4275 0.4650 0.5025 0.8250 ;
        RECT 0.3825 0.4650 0.4275 0.5850 ;
        RECT 0.2625 0.2475 0.3675 0.3900 ;
        RECT 0.3075 0.6600 0.3525 0.8250 ;
        RECT 0.2325 0.4800 0.3075 0.8250 ;
        RECT 0.1500 0.4800 0.2325 0.5550 ;
        LAYER VIA1 ;
        RECT 1.7925 0.3900 1.8675 0.4650 ;
        RECT 1.5375 0.8100 1.6125 0.8850 ;
        LAYER M2 ;
        RECT 1.8525 0.3525 1.8825 0.5025 ;
        RECT 1.7775 0.3525 1.8525 0.8700 ;
        RECT 1.6500 0.7950 1.7775 0.8700 ;
        RECT 1.5000 0.7950 1.6500 0.9000 ;
    END
END OR4_0111


MACRO OR4_1000
    CLASS CORE ;
    FOREIGN OR4_1000 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.2600 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 1.1475 0.1500 1.2225 0.9000 ;
        RECT 1.0950 0.1500 1.1475 0.3825 ;
        RECT 1.0950 0.6675 1.1475 0.9000 ;
        END
    END Z
    PIN A4
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.1425 0.4650 0.2400 0.5850 ;
        RECT 0.0675 0.3675 0.1425 0.6825 ;
        END
    END A4
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.4275 0.8625 0.8925 0.9375 ;
        RECT 0.3525 0.5550 0.4275 0.9375 ;
        VIA 0.3900 0.6675 VIA12_square ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.6600 0.7125 1.1250 0.7875 ;
        RECT 0.5100 0.6225 0.6600 0.7875 ;
        VIA 0.5850 0.6750 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.7575 0.2625 0.8325 0.5925 ;
        RECT 0.2925 0.2625 0.7575 0.3375 ;
        VIA 0.7950 0.4800 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.0050 -0.0750 1.2600 0.0750 ;
        RECT 0.8850 -0.0750 1.0050 0.1800 ;
        RECT 0.5850 -0.0750 0.8850 0.0750 ;
        RECT 0.4650 -0.0750 0.5850 0.1800 ;
        RECT 0.1650 -0.0750 0.4650 0.0750 ;
        RECT 0.0450 -0.0750 0.1650 0.2475 ;
        RECT 0.0000 -0.0750 0.0450 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.0050 0.9750 1.2600 1.1250 ;
        RECT 0.8850 0.8700 1.0050 1.1250 ;
        RECT 0.0000 0.9750 0.8850 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.1250 0.1575 1.1850 0.2175 ;
        RECT 1.1250 0.8175 1.1850 0.8775 ;
        RECT 1.0125 0.4950 1.0725 0.5550 ;
        RECT 0.9150 0.1200 0.9750 0.1800 ;
        RECT 0.9150 0.8700 0.9750 0.9300 ;
        RECT 0.8100 0.4875 0.8700 0.5475 ;
        RECT 0.7050 0.1725 0.7650 0.2325 ;
        RECT 0.5925 0.4875 0.6525 0.5475 ;
        RECT 0.4950 0.1200 0.5550 0.1800 ;
        RECT 0.3825 0.4800 0.4425 0.5400 ;
        RECT 0.2850 0.1800 0.3450 0.2400 ;
        RECT 0.1800 0.4950 0.2400 0.5550 ;
        RECT 0.0750 0.1575 0.1350 0.2175 ;
        RECT 0.0750 0.8325 0.1350 0.8925 ;
        LAYER M1 ;
        RECT 1.0200 0.4650 1.0725 0.5850 ;
        RECT 0.9450 0.2550 1.0200 0.7950 ;
        RECT 0.7875 0.2550 0.9450 0.3300 ;
        RECT 0.8100 0.7200 0.9450 0.7950 ;
        RECT 0.7275 0.4050 0.8700 0.6450 ;
        RECT 0.7350 0.7200 0.8100 0.9000 ;
        RECT 0.6825 0.1500 0.7875 0.3300 ;
        RECT 0.1500 0.8250 0.7350 0.9000 ;
        RECT 0.3675 0.2550 0.6825 0.3300 ;
        RECT 0.5175 0.4050 0.6525 0.7500 ;
        RECT 0.3300 0.4050 0.4425 0.7500 ;
        RECT 0.2625 0.1575 0.3675 0.3300 ;
        RECT 0.0450 0.7950 0.1500 0.9000 ;
    END
END OR4_1000


MACRO OR4_1010
    CLASS CORE ;
    FOREIGN OR4_1010 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.2600 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 1.1475 0.2175 1.2225 0.8325 ;
        RECT 1.1250 0.2175 1.1475 0.3825 ;
        RECT 1.1175 0.6675 1.1475 0.8325 ;
        END
    END Z
    PIN A4
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.2175 0.4500 0.2925 0.8325 ;
        RECT 0.1875 0.4500 0.2175 0.5700 ;
        END
    END A4
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.3900 0.4425 0.4950 0.8325 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.5700 0.4500 0.6600 0.8325 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.8250 0.4050 0.9000 0.5475 ;
        RECT 0.7350 0.4050 0.8250 0.8325 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.0050 -0.0750 1.2600 0.0750 ;
        RECT 0.8850 -0.0750 1.0050 0.1800 ;
        RECT 0.5850 -0.0750 0.8850 0.0750 ;
        RECT 0.4650 -0.0750 0.5850 0.1800 ;
        RECT 0.1650 -0.0750 0.4650 0.0750 ;
        RECT 0.0450 -0.0750 0.1650 0.2175 ;
        RECT 0.0000 -0.0750 0.0450 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.0125 0.9750 1.2600 1.1250 ;
        RECT 0.9075 0.6675 1.0125 1.1250 ;
        RECT 0.0000 0.9750 0.9075 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.1250 0.2700 1.1850 0.3300 ;
        RECT 1.1250 0.7200 1.1850 0.7800 ;
        RECT 1.0125 0.4725 1.0725 0.5325 ;
        RECT 0.9150 0.1200 0.9750 0.1800 ;
        RECT 0.9150 0.6975 0.9750 0.7575 ;
        RECT 0.9150 0.8625 0.9750 0.9225 ;
        RECT 0.8100 0.4650 0.8700 0.5250 ;
        RECT 0.7050 0.1725 0.7650 0.2325 ;
        RECT 0.5925 0.4875 0.6525 0.5475 ;
        RECT 0.4950 0.1200 0.5550 0.1800 ;
        RECT 0.3900 0.4800 0.4500 0.5400 ;
        RECT 0.2850 0.1800 0.3450 0.2400 ;
        RECT 0.1875 0.4800 0.2475 0.5400 ;
        RECT 0.0750 0.1575 0.1350 0.2175 ;
        RECT 0.0750 0.7500 0.1350 0.8100 ;
        LAYER M1 ;
        RECT 1.0500 0.4425 1.0725 0.5625 ;
        RECT 0.9750 0.2550 1.0500 0.5625 ;
        RECT 0.7875 0.2550 0.9750 0.3300 ;
        RECT 0.6825 0.1500 0.7875 0.3300 ;
        RECT 0.3675 0.2550 0.6825 0.3300 ;
        RECT 0.2625 0.1575 0.3675 0.3675 ;
        RECT 0.1125 0.2925 0.2625 0.3675 ;
        RECT 0.1125 0.7200 0.1425 0.8400 ;
        RECT 0.0375 0.2925 0.1125 0.8400 ;
    END
END OR4_1010


VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
  MACRO PLL_1011
    CLASS BLOCK ;
    FOREIGN PLL_1011 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 181.9500 BY 183.6600 ;
    SYMMETRY X Y ;
  PIN BWADJ_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 111.7200 0.0000 111.8250 0.0750 ;
    END
  END BWADJ_0
  PIN BWADJ_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 112.5000 0.0000 112.6050 0.0750 ;
    END
  END BWADJ_1
  PIN BWADJ_2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 113.2800 0.0000 113.3850 0.0750 ;
    END
  END BWADJ_2
  PIN BWADJ_3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 114.0600 0.0000 114.1650 0.0750 ;
    END
  END BWADJ_3
  PIN BWADJ_4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 114.8400 0.0000 114.9450 0.0750 ;
    END
  END BWADJ_4
  PIN BWADJ_5
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 115.6200 0.0000 115.7250 0.0750 ;
    END
  END BWADJ_5
  PIN BYPASS
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 110.3550 0.0000 110.4600 0.0750 ;
    END
  END BYPASS
  PIN CLKF_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 145.0650 0.0000 145.1700 0.0750 ;
    END
  END CLKF_0
  PIN CLKF_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 144.6750 0.0000 144.7800 0.0750 ;
    END
  END CLKF_1
  PIN CLKF_2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 144.2850 0.0000 144.3900 0.0750 ;
    END
  END CLKF_2
  PIN CLKF_3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 154.8150 0.0000 154.9200 0.0750 ;
    END
  END CLKF_3
  PIN CLKF_4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 154.0350 0.0000 154.1400 0.0750 ;
    END
  END CLKF_4
  PIN CLKF_5
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 153.2550 0.0000 153.3600 0.0750 ;
    END
  END CLKF_5
  PIN CLKOD_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 140.3850 0.0000 140.4900 0.0750 ;
    END
  END CLKOD_0
  PIN CLKOD_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 154.4250 0.0000 154.5300 0.0750 ;
    END
  END CLKOD_1
  PIN CLKOD_2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 152.8650 0.0000 152.9700 0.0750 ;
    END
  END CLKOD_2
  PIN CLKOD_3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 153.6450 0.0000 153.7500 0.0750 ;
    END
  END CLKOD_3
  PIN CLKOUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 134.8425 0.0000 135.1125 0.0750 ;
    END
  END CLKOUT
  PIN CLKR_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 111.1350 0.0000 111.2400 0.0750 ;
    END
  END CLKR_0
  PIN CLKR_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 124.0050 0.0000 124.1100 0.0750 ;
    END
  END CLKR_1
  PIN CLKR_2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 125.1750 0.0000 125.2800 0.0750 ;
    END
  END CLKR_2
  PIN CLKR_3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 125.5650 0.0000 125.6700 0.0750 ;
    END
  END CLKR_3
  PIN FBSLIP
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 120.0900 0.0000 120.2250 0.0750 ;
    END
  END FBSLIP
  PIN FCLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 127.5150 0.0000 127.6200 0.0750 ;
    END
  END FCLK
  PIN INTFB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 128.2950 0.0000 128.4000 0.0750 ;
    END
  END INTFB
  PIN PWRDN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 118.1550 0.0000 118.2600 0.0750 ;
    END
  END PWRDN
  PIN RCLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 125.9550 0.0000 126.0600 0.0750 ;
    END
  END RCLK
  PIN RESET
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 109.9650 0.0000 110.0700 0.0750 ;
    END
  END RESET
  PIN RFSLIP
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 119.7000 0.0000 119.8350 0.0750 ;
    END
  END RFSLIP
  PIN TEST
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 126.7350 0.0000 126.8400 0.0750 ;
    END
  END TEST
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M6 ;
        RECT 105.1200 0.0000 106.7700 0.0750 ;
      LAYER M6 ;
        RECT 129.8700 0.0000 131.5200 0.0750 ;
      LAYER M6 ;
        RECT 135.8850 0.0000 137.5350 0.0750 ;
      LAYER M6 ;
        RECT 147.1950 0.0000 148.8450 0.0750 ;
    END
  END VDD
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M4 ;
        RECT 0.0000 23.7000 0.0750 26.3250 ;
      LAYER M4 ;
        RECT 0.0000 31.9500 0.0750 34.5750 ;
      LAYER M4 ;
        RECT 0.0000 40.2000 0.0750 42.8250 ;
      LAYER M4 ;
        RECT 0.0000 48.4500 0.0750 51.0750 ;
      LAYER M4 ;
        RECT 0.0000 56.7000 0.0750 59.3250 ;
      LAYER M4 ;
        RECT 0.0000 64.9500 0.0750 67.5750 ;
      LAYER M4 ;
        RECT 0.0000 73.2000 0.0750 75.8250 ;
      LAYER M4 ;
        RECT 0.0000 81.4500 0.0750 84.0750 ;
    END
  END VDDA
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M6 ;
        RECT 107.5950 0.0000 109.2450 0.0750 ;
      LAYER M6 ;
        RECT 132.3450 0.0000 133.9950 0.0750 ;
      LAYER M6 ;
        RECT 138.3600 0.0000 140.0100 0.0750 ;
      LAYER M6 ;
        RECT 149.6700 0.0000 151.3200 0.0750 ;
    END
  END VSS
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M4 ;
        RECT 0.0000 27.8250 0.0750 30.4500 ;
      LAYER M4 ;
        RECT 0.0000 36.0750 0.0750 38.7000 ;
      LAYER M4 ;
        RECT 0.0000 44.3250 0.0750 46.9500 ;
      LAYER M4 ;
        RECT 0.0000 52.5750 0.0750 55.2000 ;
      LAYER M4 ;
        RECT 0.0000 60.8250 0.0750 63.4500 ;
      LAYER M4 ;
        RECT 0.0000 69.0750 0.0750 71.7000 ;
      LAYER M4 ;
        RECT 0.0000 77.3250 0.0750 79.9500 ;
      LAYER M4 ;
        RECT 0.0000 85.5750 0.0750 88.2000 ;
    END
  END VSSA
  OBS
    LAYER M1 ;
        RECT 0.2100 0.2100 181.7400 183.4500 ;
    LAYER M2 ;
        RECT 0.2100 0.2100 181.7400 183.4500 ;
    LAYER M3 ;
        RECT 0.2100 0.2100 181.7400 183.4500 ;
    LAYER M4 ;
        RECT 0.2100 0.2100 181.7400 183.4500 ;
    LAYER M5 ;
        RECT 0.2100 0.2100 181.7400 183.4500 ;
    LAYER M6 ;
        RECT 0.2100 0.2100 181.7400 183.4500 ;
  END
END PLL_1011


VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO SRAM2048x32M4_1001
	CLASS BLOCK ;
	FOREIGN SRAM2048x32M4_1001 0.0 0.0 ;
	ORIGIN 0.0 0.0 ;
    SIZE 242.7075 BY 141.6150 ;
	SYMMETRY X Y ;
	PIN AM[0]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
        RECT 242.4375 58.0950 242.7075 58.3200 ;
			LAYER M2 ;
        RECT 242.4375 58.0950 242.7075 58.3200 ;
			LAYER M3 ;
        RECT 242.4375 58.0950 242.7075 58.3200 ;
		END
	END AM[0]
	PIN AM[10]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
        RECT 242.4375 63.4050 242.7075 63.6300 ;
			LAYER M2 ;
        RECT 242.4375 63.4050 242.7075 63.6300 ;
			LAYER M1 ;
        RECT 242.4375 63.4050 242.7075 63.6300 ;
		END
	END AM[10]
	PIN AM[1]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
        RECT 242.4375 59.5800 242.7075 59.8050 ;
			LAYER M1 ;
        RECT 242.4375 59.5800 242.7075 59.8050 ;
			LAYER M3 ;
        RECT 242.4375 59.5800 242.7075 59.8050 ;
		END
	END AM[1]
	PIN AM[2]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
        RECT 242.4375 70.9500 242.7075 71.1750 ;
			LAYER M2 ;
        RECT 242.4375 70.9500 242.7075 71.1750 ;
			LAYER M1 ;
        RECT 242.4375 70.9500 242.7075 71.1750 ;
		END
	END AM[2]
	PIN AM[3]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
        RECT 242.4375 71.9100 242.7075 72.1350 ;
			LAYER M2 ;
        RECT 242.4375 71.9100 242.7075 72.1350 ;
			LAYER M1 ;
        RECT 242.4375 71.9100 242.7075 72.1350 ;
		END
	END AM[3]
	PIN AM[4]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
        RECT 242.4375 73.7850 242.7075 74.0100 ;
			LAYER M1 ;
        RECT 242.4375 73.7850 242.7075 74.0100 ;
			LAYER M3 ;
        RECT 242.4375 73.7850 242.7075 74.0100 ;
		END
	END AM[4]
	PIN AM[5]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
        RECT 242.4375 69.0750 242.7075 69.3000 ;
			LAYER M2 ;
        RECT 242.4375 69.0750 242.7075 69.3000 ;
			LAYER M1 ;
        RECT 242.4375 69.0750 242.7075 69.3000 ;
		END
	END AM[5]
	PIN AM[6]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
        RECT 242.4375 68.1150 242.7075 68.3400 ;
			LAYER M1 ;
        RECT 242.4375 68.1150 242.7075 68.3400 ;
			LAYER M2 ;
        RECT 242.4375 68.1150 242.7075 68.3400 ;
		END
	END AM[6]
	PIN AM[7]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
        RECT 242.4375 66.2400 242.7075 66.4650 ;
			LAYER M3 ;
        RECT 242.4375 66.2400 242.7075 66.4650 ;
			LAYER M2 ;
        RECT 242.4375 66.2400 242.7075 66.4650 ;
		END
	END AM[7]
	PIN AM[8]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
        RECT 242.4375 60.5700 242.7075 60.7950 ;
			LAYER M3 ;
        RECT 242.4375 60.5700 242.7075 60.7950 ;
			LAYER M2 ;
        RECT 242.4375 60.5700 242.7075 60.7950 ;
		END
	END AM[8]
	PIN AM[9]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
        RECT 242.4375 62.4450 242.7075 62.6700 ;
			LAYER M1 ;
        RECT 242.4375 62.4450 242.7075 62.6700 ;
			LAYER M3 ;
        RECT 242.4375 62.4450 242.7075 62.6700 ;
		END
	END AM[9]
	PIN A[0]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
        RECT 242.4375 58.5900 242.7075 58.8150 ;
			LAYER M2 ;
        RECT 242.4375 58.5900 242.7075 58.8150 ;
			LAYER M1 ;
        RECT 242.4375 58.5900 242.7075 58.8150 ;
		END
	END A[0]
	PIN A[10]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
        RECT 242.4375 64.0950 242.7075 64.3200 ;
			LAYER M2 ;
        RECT 242.4375 64.0950 242.7075 64.3200 ;
			LAYER M1 ;
        RECT 242.4375 64.0950 242.7075 64.3200 ;
		END
	END A[10]
	PIN A[1]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
        RECT 242.4375 59.0850 242.7075 59.3100 ;
			LAYER M2 ;
        RECT 242.4375 59.0850 242.7075 59.3100 ;
			LAYER M1 ;
        RECT 242.4375 59.0850 242.7075 59.3100 ;
		END
	END A[1]
	PIN A[2]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
        RECT 242.4375 70.2600 242.7075 70.4850 ;
			LAYER M2 ;
        RECT 242.4375 70.2600 242.7075 70.4850 ;
			LAYER M1 ;
        RECT 242.4375 70.2600 242.7075 70.4850 ;
		END
	END A[2]
	PIN A[3]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
        RECT 242.4375 72.6000 242.7075 72.8250 ;
			LAYER M2 ;
        RECT 242.4375 72.6000 242.7075 72.8250 ;
			LAYER M3 ;
        RECT 242.4375 72.6000 242.7075 72.8250 ;
		END
	END A[3]
	PIN A[4]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
        RECT 242.4375 73.0950 242.7075 73.3200 ;
			LAYER M2 ;
        RECT 242.4375 73.0950 242.7075 73.3200 ;
			LAYER M3 ;
        RECT 242.4375 73.0950 242.7075 73.3200 ;
		END
	END A[4]
	PIN A[5]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
        RECT 242.4375 69.7650 242.7075 69.9900 ;
			LAYER M1 ;
        RECT 242.4375 69.7650 242.7075 69.9900 ;
			LAYER M2 ;
        RECT 242.4375 69.7650 242.7075 69.9900 ;
		END
	END A[5]
	PIN A[6]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
        RECT 242.4375 67.4250 242.7075 67.6500 ;
			LAYER M1 ;
        RECT 242.4375 67.4250 242.7075 67.6500 ;
			LAYER M3 ;
        RECT 242.4375 67.4250 242.7075 67.6500 ;
		END
	END A[6]
	PIN A[7]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
        RECT 242.4375 66.9300 242.7075 67.1550 ;
			LAYER M2 ;
        RECT 242.4375 66.9300 242.7075 67.1550 ;
			LAYER M1 ;
        RECT 242.4375 66.9300 242.7075 67.1550 ;
		END
	END A[7]
	PIN A[8]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
        RECT 242.4375 61.2600 242.7075 61.4850 ;
			LAYER M3 ;
        RECT 242.4375 61.2600 242.7075 61.4850 ;
			LAYER M1 ;
        RECT 242.4375 61.2600 242.7075 61.4850 ;
		END
	END A[8]
	PIN A[9]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
        RECT 242.4375 61.7550 242.7075 61.9800 ;
			LAYER M3 ;
        RECT 242.4375 61.7550 242.7075 61.9800 ;
			LAYER M1 ;
        RECT 242.4375 61.7550 242.7075 61.9800 ;
		END
	END A[9]
	PIN BIST
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
        RECT 242.4375 77.5275 242.7075 77.7525 ;
			LAYER M3 ;
        RECT 242.4375 77.5275 242.7075 77.7525 ;
			LAYER M2 ;
        RECT 242.4375 77.5275 242.7075 77.7525 ;
		END
	END BIST
	PIN BWEBM[0]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
        RECT 242.4375 1.4025 242.7075 1.6275 ;
			LAYER M2 ;
        RECT 242.4375 1.4025 242.7075 1.6275 ;
			LAYER M1 ;
        RECT 242.4375 1.4025 242.7075 1.6275 ;
		END
	END BWEBM[0]
	PIN BWEBM[10]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
        RECT 242.4375 36.2025 242.7075 36.4275 ;
			LAYER M2 ;
        RECT 242.4375 36.2025 242.7075 36.4275 ;
			LAYER M3 ;
        RECT 242.4375 36.2025 242.7075 36.4275 ;
		END
	END BWEBM[10]
	PIN BWEBM[11]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
        RECT 242.4375 39.6825 242.7075 39.9075 ;
			LAYER M2 ;
        RECT 242.4375 39.6825 242.7075 39.9075 ;
			LAYER M1 ;
        RECT 242.4375 39.6825 242.7075 39.9075 ;
		END
	END BWEBM[11]
	PIN BWEBM[12]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
        RECT 242.4375 43.1625 242.7075 43.3875 ;
			LAYER M3 ;
        RECT 242.4375 43.1625 242.7075 43.3875 ;
			LAYER M1 ;
        RECT 242.4375 43.1625 242.7075 43.3875 ;
		END
	END BWEBM[12]
	PIN BWEBM[13]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
        RECT 242.4375 46.6425 242.7075 46.8675 ;
			LAYER M2 ;
        RECT 242.4375 46.6425 242.7075 46.8675 ;
			LAYER M3 ;
        RECT 242.4375 46.6425 242.7075 46.8675 ;
		END
	END BWEBM[13]
	PIN BWEBM[14]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
        RECT 242.4375 50.1225 242.7075 50.3475 ;
			LAYER M1 ;
        RECT 242.4375 50.1225 242.7075 50.3475 ;
			LAYER M3 ;
        RECT 242.4375 50.1225 242.7075 50.3475 ;
		END
	END BWEBM[14]
	PIN BWEBM[15]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
        RECT 242.4375 53.6025 242.7075 53.8275 ;
			LAYER M1 ;
        RECT 242.4375 53.6025 242.7075 53.8275 ;
			LAYER M3 ;
        RECT 242.4375 53.6025 242.7075 53.8275 ;
		END
	END BWEBM[15]
	PIN BWEBM[16]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
        RECT 242.4375 84.8325 242.7075 85.0575 ;
			LAYER M2 ;
        RECT 242.4375 84.8325 242.7075 85.0575 ;
			LAYER M1 ;
        RECT 242.4375 84.8325 242.7075 85.0575 ;
		END
	END BWEBM[16]
	PIN BWEBM[17]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
        RECT 242.4375 88.3125 242.7075 88.5375 ;
			LAYER M3 ;
        RECT 242.4375 88.3125 242.7075 88.5375 ;
			LAYER M1 ;
        RECT 242.4375 88.3125 242.7075 88.5375 ;
		END
	END BWEBM[17]
	PIN BWEBM[18]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
        RECT 242.4375 91.7925 242.7075 92.0175 ;
			LAYER M2 ;
        RECT 242.4375 91.7925 242.7075 92.0175 ;
			LAYER M3 ;
        RECT 242.4375 91.7925 242.7075 92.0175 ;
		END
	END BWEBM[18]
	PIN BWEBM[19]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
        RECT 242.4375 95.2725 242.7075 95.4975 ;
			LAYER M1 ;
        RECT 242.4375 95.2725 242.7075 95.4975 ;
			LAYER M2 ;
        RECT 242.4375 95.2725 242.7075 95.4975 ;
		END
	END BWEBM[19]
	PIN BWEBM[1]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
        RECT 242.4375 4.8825 242.7075 5.1075 ;
			LAYER M2 ;
        RECT 242.4375 4.8825 242.7075 5.1075 ;
			LAYER M1 ;
        RECT 242.4375 4.8825 242.7075 5.1075 ;
		END
	END BWEBM[1]
	PIN BWEBM[20]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
        RECT 242.4375 98.7525 242.7075 98.9775 ;
			LAYER M3 ;
        RECT 242.4375 98.7525 242.7075 98.9775 ;
			LAYER M2 ;
        RECT 242.4375 98.7525 242.7075 98.9775 ;
		END
	END BWEBM[20]
	PIN BWEBM[21]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
        RECT 242.4375 102.2325 242.7075 102.4575 ;
			LAYER M1 ;
        RECT 242.4375 102.2325 242.7075 102.4575 ;
			LAYER M3 ;
        RECT 242.4375 102.2325 242.7075 102.4575 ;
		END
	END BWEBM[21]
	PIN BWEBM[22]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
        RECT 242.4375 105.7125 242.7075 105.9375 ;
			LAYER M1 ;
        RECT 242.4375 105.7125 242.7075 105.9375 ;
			LAYER M2 ;
        RECT 242.4375 105.7125 242.7075 105.9375 ;
		END
	END BWEBM[22]
	PIN BWEBM[23]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
        RECT 242.4375 109.1925 242.7075 109.4175 ;
			LAYER M3 ;
        RECT 242.4375 109.1925 242.7075 109.4175 ;
			LAYER M2 ;
        RECT 242.4375 109.1925 242.7075 109.4175 ;
		END
	END BWEBM[23]
	PIN BWEBM[24]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
        RECT 242.4375 112.6725 242.7075 112.8975 ;
			LAYER M1 ;
        RECT 242.4375 112.6725 242.7075 112.8975 ;
			LAYER M2 ;
        RECT 242.4375 112.6725 242.7075 112.8975 ;
		END
	END BWEBM[24]
	PIN BWEBM[25]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
        RECT 242.4375 116.1525 242.7075 116.3775 ;
			LAYER M2 ;
        RECT 242.4375 116.1525 242.7075 116.3775 ;
			LAYER M3 ;
        RECT 242.4375 116.1525 242.7075 116.3775 ;
		END
	END BWEBM[25]
	PIN BWEBM[26]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
        RECT 242.4375 119.6325 242.7075 119.8575 ;
			LAYER M2 ;
        RECT 242.4375 119.6325 242.7075 119.8575 ;
			LAYER M3 ;
        RECT 242.4375 119.6325 242.7075 119.8575 ;
		END
	END BWEBM[26]
	PIN BWEBM[27]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
        RECT 242.4375 123.1125 242.7075 123.3375 ;
			LAYER M2 ;
        RECT 242.4375 123.1125 242.7075 123.3375 ;
			LAYER M3 ;
        RECT 242.4375 123.1125 242.7075 123.3375 ;
		END
	END BWEBM[27]
	PIN BWEBM[28]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
        RECT 242.4375 126.5925 242.7075 126.8175 ;
			LAYER M1 ;
        RECT 242.4375 126.5925 242.7075 126.8175 ;
			LAYER M2 ;
        RECT 242.4375 126.5925 242.7075 126.8175 ;
		END
	END BWEBM[28]
	PIN BWEBM[29]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
        RECT 242.4375 130.0725 242.7075 130.2975 ;
			LAYER M3 ;
        RECT 242.4375 130.0725 242.7075 130.2975 ;
			LAYER M1 ;
        RECT 242.4375 130.0725 242.7075 130.2975 ;
		END
	END BWEBM[29]
	PIN BWEBM[2]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
        RECT 242.4375 8.3625 242.7075 8.5875 ;
			LAYER M2 ;
        RECT 242.4375 8.3625 242.7075 8.5875 ;
			LAYER M3 ;
        RECT 242.4375 8.3625 242.7075 8.5875 ;
		END
	END BWEBM[2]
	PIN BWEBM[30]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
        RECT 242.4375 133.5525 242.7075 133.7775 ;
			LAYER M1 ;
        RECT 242.4375 133.5525 242.7075 133.7775 ;
			LAYER M2 ;
        RECT 242.4375 133.5525 242.7075 133.7775 ;
		END
	END BWEBM[30]
	PIN BWEBM[31]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
        RECT 242.4375 137.0325 242.7075 137.2575 ;
			LAYER M1 ;
        RECT 242.4375 137.0325 242.7075 137.2575 ;
			LAYER M3 ;
        RECT 242.4375 137.0325 242.7075 137.2575 ;
		END
	END BWEBM[31]
	PIN BWEBM[3]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
        RECT 242.4375 11.8425 242.7075 12.0675 ;
			LAYER M3 ;
        RECT 242.4375 11.8425 242.7075 12.0675 ;
			LAYER M1 ;
        RECT 242.4375 11.8425 242.7075 12.0675 ;
		END
	END BWEBM[3]
	PIN BWEBM[4]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
        RECT 242.4375 15.3225 242.7075 15.5475 ;
			LAYER M3 ;
        RECT 242.4375 15.3225 242.7075 15.5475 ;
			LAYER M2 ;
        RECT 242.4375 15.3225 242.7075 15.5475 ;
		END
	END BWEBM[4]
	PIN BWEBM[5]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
        RECT 242.4375 18.8025 242.7075 19.0275 ;
			LAYER M3 ;
        RECT 242.4375 18.8025 242.7075 19.0275 ;
			LAYER M1 ;
        RECT 242.4375 18.8025 242.7075 19.0275 ;
		END
	END BWEBM[5]
	PIN BWEBM[6]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
        RECT 242.4375 22.2825 242.7075 22.5075 ;
			LAYER M1 ;
        RECT 242.4375 22.2825 242.7075 22.5075 ;
			LAYER M2 ;
        RECT 242.4375 22.2825 242.7075 22.5075 ;
		END
	END BWEBM[6]
	PIN BWEBM[7]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
        RECT 242.4375 25.7625 242.7075 25.9875 ;
			LAYER M1 ;
        RECT 242.4375 25.7625 242.7075 25.9875 ;
			LAYER M2 ;
        RECT 242.4375 25.7625 242.7075 25.9875 ;
		END
	END BWEBM[7]
	PIN BWEBM[8]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
        RECT 242.4375 29.2425 242.7075 29.4675 ;
			LAYER M3 ;
        RECT 242.4375 29.2425 242.7075 29.4675 ;
			LAYER M1 ;
        RECT 242.4375 29.2425 242.7075 29.4675 ;
		END
	END BWEBM[8]
	PIN BWEBM[9]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
        RECT 242.4375 32.7225 242.7075 32.9475 ;
			LAYER M3 ;
        RECT 242.4375 32.7225 242.7075 32.9475 ;
			LAYER M2 ;
        RECT 242.4375 32.7225 242.7075 32.9475 ;
		END
	END BWEBM[9]
	PIN BWEB[0]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
        RECT 242.4375 1.8975 242.7075 2.1225 ;
			LAYER M2 ;
        RECT 242.4375 1.8975 242.7075 2.1225 ;
			LAYER M1 ;
        RECT 242.4375 1.8975 242.7075 2.1225 ;
		END
	END BWEB[0]
	PIN BWEB[10]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
        RECT 242.4375 36.6975 242.7075 36.9225 ;
			LAYER M1 ;
        RECT 242.4375 36.6975 242.7075 36.9225 ;
			LAYER M2 ;
        RECT 242.4375 36.6975 242.7075 36.9225 ;
		END
	END BWEB[10]
	PIN BWEB[11]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
        RECT 242.4375 40.1775 242.7075 40.4025 ;
			LAYER M1 ;
        RECT 242.4375 40.1775 242.7075 40.4025 ;
			LAYER M3 ;
        RECT 242.4375 40.1775 242.7075 40.4025 ;
		END
	END BWEB[11]
	PIN BWEB[12]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
        RECT 242.4375 43.6575 242.7075 43.8825 ;
			LAYER M3 ;
        RECT 242.4375 43.6575 242.7075 43.8825 ;
			LAYER M1 ;
        RECT 242.4375 43.6575 242.7075 43.8825 ;
		END
	END BWEB[12]
	PIN BWEB[13]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
        RECT 242.4375 47.1375 242.7075 47.3625 ;
			LAYER M3 ;
        RECT 242.4375 47.1375 242.7075 47.3625 ;
			LAYER M1 ;
        RECT 242.4375 47.1375 242.7075 47.3625 ;
		END
	END BWEB[13]
	PIN BWEB[14]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
        RECT 242.4375 50.6175 242.7075 50.8425 ;
			LAYER M1 ;
        RECT 242.4375 50.6175 242.7075 50.8425 ;
			LAYER M3 ;
        RECT 242.4375 50.6175 242.7075 50.8425 ;
		END
	END BWEB[14]
	PIN BWEB[15]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
        RECT 242.4375 54.0975 242.7075 54.3225 ;
			LAYER M2 ;
        RECT 242.4375 54.0975 242.7075 54.3225 ;
			LAYER M1 ;
        RECT 242.4375 54.0975 242.7075 54.3225 ;
		END
	END BWEB[15]
	PIN BWEB[16]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
        RECT 242.4375 85.3275 242.7075 85.5525 ;
			LAYER M3 ;
        RECT 242.4375 85.3275 242.7075 85.5525 ;
			LAYER M1 ;
        RECT 242.4375 85.3275 242.7075 85.5525 ;
		END
	END BWEB[16]
	PIN BWEB[17]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
        RECT 242.4375 88.8075 242.7075 89.0325 ;
			LAYER M1 ;
        RECT 242.4375 88.8075 242.7075 89.0325 ;
			LAYER M3 ;
        RECT 242.4375 88.8075 242.7075 89.0325 ;
		END
	END BWEB[17]
	PIN BWEB[18]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
        RECT 242.4375 92.2875 242.7075 92.5125 ;
			LAYER M3 ;
        RECT 242.4375 92.2875 242.7075 92.5125 ;
			LAYER M1 ;
        RECT 242.4375 92.2875 242.7075 92.5125 ;
		END
	END BWEB[18]
	PIN BWEB[19]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
        RECT 242.4375 95.7675 242.7075 95.9925 ;
			LAYER M2 ;
        RECT 242.4375 95.7675 242.7075 95.9925 ;
			LAYER M1 ;
        RECT 242.4375 95.7675 242.7075 95.9925 ;
		END
	END BWEB[19]
	PIN BWEB[1]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
        RECT 242.4375 5.3775 242.7075 5.6025 ;
			LAYER M2 ;
        RECT 242.4375 5.3775 242.7075 5.6025 ;
			LAYER M1 ;
        RECT 242.4375 5.3775 242.7075 5.6025 ;
		END
	END BWEB[1]
	PIN BWEB[20]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
        RECT 242.4375 99.2475 242.7075 99.4725 ;
			LAYER M3 ;
        RECT 242.4375 99.2475 242.7075 99.4725 ;
			LAYER M1 ;
        RECT 242.4375 99.2475 242.7075 99.4725 ;
		END
	END BWEB[20]
	PIN BWEB[21]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
        RECT 242.4375 102.7275 242.7075 102.9525 ;
			LAYER M3 ;
        RECT 242.4375 102.7275 242.7075 102.9525 ;
			LAYER M1 ;
        RECT 242.4375 102.7275 242.7075 102.9525 ;
		END
	END BWEB[21]
	PIN BWEB[22]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
        RECT 242.4375 106.2075 242.7075 106.4325 ;
			LAYER M3 ;
        RECT 242.4375 106.2075 242.7075 106.4325 ;
			LAYER M2 ;
        RECT 242.4375 106.2075 242.7075 106.4325 ;
		END
	END BWEB[22]
	PIN BWEB[23]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
        RECT 242.4375 109.6875 242.7075 109.9125 ;
			LAYER M2 ;
        RECT 242.4375 109.6875 242.7075 109.9125 ;
			LAYER M1 ;
        RECT 242.4375 109.6875 242.7075 109.9125 ;
		END
	END BWEB[23]
	PIN BWEB[24]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
        RECT 242.4375 113.1675 242.7075 113.3925 ;
			LAYER M1 ;
        RECT 242.4375 113.1675 242.7075 113.3925 ;
			LAYER M3 ;
        RECT 242.4375 113.1675 242.7075 113.3925 ;
		END
	END BWEB[24]
	PIN BWEB[25]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
        RECT 242.4375 116.6475 242.7075 116.8725 ;
			LAYER M2 ;
        RECT 242.4375 116.6475 242.7075 116.8725 ;
			LAYER M3 ;
        RECT 242.4375 116.6475 242.7075 116.8725 ;
		END
	END BWEB[25]
	PIN BWEB[26]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
        RECT 242.4375 120.1275 242.7075 120.3525 ;
			LAYER M1 ;
        RECT 242.4375 120.1275 242.7075 120.3525 ;
			LAYER M3 ;
        RECT 242.4375 120.1275 242.7075 120.3525 ;
		END
	END BWEB[26]
	PIN BWEB[27]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
        RECT 242.4375 123.6075 242.7075 123.8325 ;
			LAYER M3 ;
        RECT 242.4375 123.6075 242.7075 123.8325 ;
			LAYER M2 ;
        RECT 242.4375 123.6075 242.7075 123.8325 ;
		END
	END BWEB[27]
	PIN BWEB[28]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
        RECT 242.4375 127.0875 242.7075 127.3125 ;
			LAYER M1 ;
        RECT 242.4375 127.0875 242.7075 127.3125 ;
			LAYER M2 ;
        RECT 242.4375 127.0875 242.7075 127.3125 ;
		END
	END BWEB[28]
	PIN BWEB[29]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
        RECT 242.4375 130.5675 242.7075 130.7925 ;
			LAYER M2 ;
        RECT 242.4375 130.5675 242.7075 130.7925 ;
			LAYER M3 ;
        RECT 242.4375 130.5675 242.7075 130.7925 ;
		END
	END BWEB[29]
	PIN BWEB[2]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
        RECT 242.4375 8.8575 242.7075 9.0825 ;
			LAYER M1 ;
        RECT 242.4375 8.8575 242.7075 9.0825 ;
			LAYER M3 ;
        RECT 242.4375 8.8575 242.7075 9.0825 ;
		END
	END BWEB[2]
	PIN BWEB[30]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
        RECT 242.4375 134.0475 242.7075 134.2725 ;
			LAYER M2 ;
        RECT 242.4375 134.0475 242.7075 134.2725 ;
			LAYER M1 ;
        RECT 242.4375 134.0475 242.7075 134.2725 ;
		END
	END BWEB[30]
	PIN BWEB[31]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
        RECT 242.4375 137.5275 242.7075 137.7525 ;
			LAYER M3 ;
        RECT 242.4375 137.5275 242.7075 137.7525 ;
			LAYER M2 ;
        RECT 242.4375 137.5275 242.7075 137.7525 ;
		END
	END BWEB[31]
	PIN BWEB[3]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
        RECT 242.4375 12.3375 242.7075 12.5625 ;
			LAYER M2 ;
        RECT 242.4375 12.3375 242.7075 12.5625 ;
			LAYER M1 ;
        RECT 242.4375 12.3375 242.7075 12.5625 ;
		END
	END BWEB[3]
	PIN BWEB[4]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
        RECT 242.4375 15.8175 242.7075 16.0425 ;
			LAYER M3 ;
        RECT 242.4375 15.8175 242.7075 16.0425 ;
			LAYER M1 ;
        RECT 242.4375 15.8175 242.7075 16.0425 ;
		END
	END BWEB[4]
	PIN BWEB[5]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
        RECT 242.4375 19.2975 242.7075 19.5225 ;
			LAYER M2 ;
        RECT 242.4375 19.2975 242.7075 19.5225 ;
			LAYER M1 ;
        RECT 242.4375 19.2975 242.7075 19.5225 ;
		END
	END BWEB[5]
	PIN BWEB[6]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
        RECT 242.4375 22.7775 242.7075 23.0025 ;
			LAYER M1 ;
        RECT 242.4375 22.7775 242.7075 23.0025 ;
			LAYER M2 ;
        RECT 242.4375 22.7775 242.7075 23.0025 ;
		END
	END BWEB[6]
	PIN BWEB[7]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
        RECT 242.4375 26.2575 242.7075 26.4825 ;
			LAYER M3 ;
        RECT 242.4375 26.2575 242.7075 26.4825 ;
			LAYER M2 ;
        RECT 242.4375 26.2575 242.7075 26.4825 ;
		END
	END BWEB[7]
	PIN BWEB[8]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
        RECT 242.4375 29.7375 242.7075 29.9625 ;
			LAYER M2 ;
        RECT 242.4375 29.7375 242.7075 29.9625 ;
			LAYER M1 ;
        RECT 242.4375 29.7375 242.7075 29.9625 ;
		END
	END BWEB[8]
	PIN BWEB[9]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
        RECT 242.4375 33.2175 242.7075 33.4425 ;
			LAYER M1 ;
        RECT 242.4375 33.2175 242.7075 33.4425 ;
			LAYER M3 ;
        RECT 242.4375 33.2175 242.7075 33.4425 ;
		END
	END BWEB[9]
	PIN CEB
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
        RECT 242.4375 75.4350 242.7075 75.6600 ;
			LAYER M3 ;
        RECT 242.4375 75.4350 242.7075 75.6600 ;
			LAYER M2 ;
        RECT 242.4375 75.4350 242.7075 75.6600 ;
		END
	END CEB
	PIN CEBM
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
        RECT 242.4375 74.7450 242.7075 74.9700 ;
			LAYER M2 ;
        RECT 242.4375 74.7450 242.7075 74.9700 ;
			LAYER M1 ;
        RECT 242.4375 74.7450 242.7075 74.9700 ;
		END
	END CEBM
	PIN CLK
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
        RECT 242.4375 80.5350 242.7075 80.7600 ;
			LAYER M1 ;
        RECT 242.4375 80.5350 242.7075 80.7600 ;
			LAYER M3 ;
        RECT 242.4375 80.5350 242.7075 80.7600 ;
		END
	END CLK
	PIN DM[0]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
        RECT 242.4375 4.3575 242.7075 4.5825 ;
			LAYER M2 ;
        RECT 242.4375 4.3575 242.7075 4.5825 ;
			LAYER M3 ;
        RECT 242.4375 4.3575 242.7075 4.5825 ;
		END
	END DM[0]
	PIN DM[10]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
        RECT 242.4375 39.1575 242.7075 39.3825 ;
			LAYER M2 ;
        RECT 242.4375 39.1575 242.7075 39.3825 ;
			LAYER M3 ;
        RECT 242.4375 39.1575 242.7075 39.3825 ;
		END
	END DM[10]
	PIN DM[11]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
        RECT 242.4375 42.6375 242.7075 42.8625 ;
			LAYER M3 ;
        RECT 242.4375 42.6375 242.7075 42.8625 ;
			LAYER M2 ;
        RECT 242.4375 42.6375 242.7075 42.8625 ;
		END
	END DM[11]
	PIN DM[12]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
        RECT 242.4375 46.1175 242.7075 46.3425 ;
			LAYER M1 ;
        RECT 242.4375 46.1175 242.7075 46.3425 ;
			LAYER M3 ;
        RECT 242.4375 46.1175 242.7075 46.3425 ;
		END
	END DM[12]
	PIN DM[13]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
        RECT 242.4375 49.5975 242.7075 49.8225 ;
			LAYER M2 ;
        RECT 242.4375 49.5975 242.7075 49.8225 ;
			LAYER M3 ;
        RECT 242.4375 49.5975 242.7075 49.8225 ;
		END
	END DM[13]
	PIN DM[14]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
        RECT 242.4375 53.0775 242.7075 53.3025 ;
			LAYER M1 ;
        RECT 242.4375 53.0775 242.7075 53.3025 ;
			LAYER M3 ;
        RECT 242.4375 53.0775 242.7075 53.3025 ;
		END
	END DM[14]
	PIN DM[15]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
        RECT 242.4375 56.5575 242.7075 56.7825 ;
			LAYER M1 ;
        RECT 242.4375 56.5575 242.7075 56.7825 ;
			LAYER M2 ;
        RECT 242.4375 56.5575 242.7075 56.7825 ;
		END
	END DM[15]
	PIN DM[16]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
        RECT 242.4375 87.7875 242.7075 88.0125 ;
			LAYER M2 ;
        RECT 242.4375 87.7875 242.7075 88.0125 ;
			LAYER M3 ;
        RECT 242.4375 87.7875 242.7075 88.0125 ;
		END
	END DM[16]
	PIN DM[17]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
        RECT 242.4375 91.2675 242.7075 91.4925 ;
			LAYER M2 ;
        RECT 242.4375 91.2675 242.7075 91.4925 ;
			LAYER M1 ;
        RECT 242.4375 91.2675 242.7075 91.4925 ;
		END
	END DM[17]
	PIN DM[18]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
        RECT 242.4375 94.7475 242.7075 94.9725 ;
			LAYER M2 ;
        RECT 242.4375 94.7475 242.7075 94.9725 ;
			LAYER M3 ;
        RECT 242.4375 94.7475 242.7075 94.9725 ;
		END
	END DM[18]
	PIN DM[19]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
        RECT 242.4375 98.2275 242.7075 98.4525 ;
			LAYER M3 ;
        RECT 242.4375 98.2275 242.7075 98.4525 ;
			LAYER M1 ;
        RECT 242.4375 98.2275 242.7075 98.4525 ;
		END
	END DM[19]
	PIN DM[1]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
        RECT 242.4375 7.8375 242.7075 8.0625 ;
			LAYER M2 ;
        RECT 242.4375 7.8375 242.7075 8.0625 ;
			LAYER M3 ;
        RECT 242.4375 7.8375 242.7075 8.0625 ;
		END
	END DM[1]
	PIN DM[20]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
        RECT 242.4375 101.7075 242.7075 101.9325 ;
			LAYER M2 ;
        RECT 242.4375 101.7075 242.7075 101.9325 ;
			LAYER M1 ;
        RECT 242.4375 101.7075 242.7075 101.9325 ;
		END
	END DM[20]
	PIN DM[21]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
        RECT 242.4375 105.1875 242.7075 105.4125 ;
			LAYER M3 ;
        RECT 242.4375 105.1875 242.7075 105.4125 ;
			LAYER M2 ;
        RECT 242.4375 105.1875 242.7075 105.4125 ;
		END
	END DM[21]
	PIN DM[22]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
        RECT 242.4375 108.6675 242.7075 108.8925 ;
			LAYER M3 ;
        RECT 242.4375 108.6675 242.7075 108.8925 ;
			LAYER M1 ;
        RECT 242.4375 108.6675 242.7075 108.8925 ;
		END
	END DM[22]
	PIN DM[23]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
        RECT 242.4375 112.1475 242.7075 112.3725 ;
			LAYER M3 ;
        RECT 242.4375 112.1475 242.7075 112.3725 ;
			LAYER M2 ;
        RECT 242.4375 112.1475 242.7075 112.3725 ;
		END
	END DM[23]
	PIN DM[24]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
        RECT 242.4375 115.6275 242.7075 115.8525 ;
			LAYER M3 ;
        RECT 242.4375 115.6275 242.7075 115.8525 ;
			LAYER M1 ;
        RECT 242.4375 115.6275 242.7075 115.8525 ;
		END
	END DM[24]
	PIN DM[25]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
        RECT 242.4375 119.1075 242.7075 119.3325 ;
			LAYER M2 ;
        RECT 242.4375 119.1075 242.7075 119.3325 ;
			LAYER M3 ;
        RECT 242.4375 119.1075 242.7075 119.3325 ;
		END
	END DM[25]
	PIN DM[26]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
        RECT 242.4375 122.5875 242.7075 122.8125 ;
			LAYER M3 ;
        RECT 242.4375 122.5875 242.7075 122.8125 ;
			LAYER M2 ;
        RECT 242.4375 122.5875 242.7075 122.8125 ;
		END
	END DM[26]
	PIN DM[27]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
        RECT 242.4375 126.0675 242.7075 126.2925 ;
			LAYER M2 ;
        RECT 242.4375 126.0675 242.7075 126.2925 ;
			LAYER M3 ;
        RECT 242.4375 126.0675 242.7075 126.2925 ;
		END
	END DM[27]
	PIN DM[28]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
        RECT 242.4375 129.5475 242.7075 129.7725 ;
			LAYER M3 ;
        RECT 242.4375 129.5475 242.7075 129.7725 ;
			LAYER M1 ;
        RECT 242.4375 129.5475 242.7075 129.7725 ;
		END
	END DM[28]
	PIN DM[29]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
        RECT 242.4375 133.0275 242.7075 133.2525 ;
			LAYER M3 ;
        RECT 242.4375 133.0275 242.7075 133.2525 ;
			LAYER M2 ;
        RECT 242.4375 133.0275 242.7075 133.2525 ;
		END
	END DM[29]
	PIN DM[2]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
        RECT 242.4375 11.3175 242.7075 11.5425 ;
			LAYER M2 ;
        RECT 242.4375 11.3175 242.7075 11.5425 ;
			LAYER M1 ;
        RECT 242.4375 11.3175 242.7075 11.5425 ;
		END
	END DM[2]
	PIN DM[30]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
        RECT 242.4375 136.5075 242.7075 136.7325 ;
			LAYER M3 ;
        RECT 242.4375 136.5075 242.7075 136.7325 ;
			LAYER M2 ;
        RECT 242.4375 136.5075 242.7075 136.7325 ;
		END
	END DM[30]
	PIN DM[31]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
        RECT 242.4375 139.9875 242.7075 140.2125 ;
			LAYER M2 ;
        RECT 242.4375 139.9875 242.7075 140.2125 ;
			LAYER M3 ;
        RECT 242.4375 139.9875 242.7075 140.2125 ;
		END
	END DM[31]
	PIN DM[3]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
        RECT 242.4375 14.7975 242.7075 15.0225 ;
			LAYER M1 ;
        RECT 242.4375 14.7975 242.7075 15.0225 ;
			LAYER M2 ;
        RECT 242.4375 14.7975 242.7075 15.0225 ;
		END
	END DM[3]
	PIN DM[4]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
        RECT 242.4375 18.2775 242.7075 18.5025 ;
			LAYER M2 ;
        RECT 242.4375 18.2775 242.7075 18.5025 ;
			LAYER M1 ;
        RECT 242.4375 18.2775 242.7075 18.5025 ;
		END
	END DM[4]
	PIN DM[5]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
        RECT 242.4375 21.7575 242.7075 21.9825 ;
			LAYER M3 ;
        RECT 242.4375 21.7575 242.7075 21.9825 ;
			LAYER M2 ;
        RECT 242.4375 21.7575 242.7075 21.9825 ;
		END
	END DM[5]
	PIN DM[6]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
        RECT 242.4375 25.2375 242.7075 25.4625 ;
			LAYER M3 ;
        RECT 242.4375 25.2375 242.7075 25.4625 ;
			LAYER M1 ;
        RECT 242.4375 25.2375 242.7075 25.4625 ;
		END
	END DM[6]
	PIN DM[7]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
        RECT 242.4375 28.7175 242.7075 28.9425 ;
			LAYER M2 ;
        RECT 242.4375 28.7175 242.7075 28.9425 ;
			LAYER M3 ;
        RECT 242.4375 28.7175 242.7075 28.9425 ;
		END
	END DM[7]
	PIN DM[8]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
        RECT 242.4375 32.1975 242.7075 32.4225 ;
			LAYER M1 ;
        RECT 242.4375 32.1975 242.7075 32.4225 ;
			LAYER M3 ;
        RECT 242.4375 32.1975 242.7075 32.4225 ;
		END
	END DM[8]
	PIN DM[9]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
        RECT 242.4375 35.6775 242.7075 35.9025 ;
			LAYER M2 ;
        RECT 242.4375 35.6775 242.7075 35.9025 ;
			LAYER M1 ;
        RECT 242.4375 35.6775 242.7075 35.9025 ;
		END
	END DM[9]
	PIN D[0]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
        RECT 242.4375 3.8625 242.7075 4.0875 ;
			LAYER M3 ;
        RECT 242.4375 3.8625 242.7075 4.0875 ;
			LAYER M2 ;
        RECT 242.4375 3.8625 242.7075 4.0875 ;
		END
	END D[0]
	PIN D[10]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
        RECT 242.4375 38.6625 242.7075 38.8875 ;
			LAYER M2 ;
        RECT 242.4375 38.6625 242.7075 38.8875 ;
			LAYER M1 ;
        RECT 242.4375 38.6625 242.7075 38.8875 ;
		END
	END D[10]
	PIN D[11]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
        RECT 242.4375 42.1425 242.7075 42.3675 ;
			LAYER M2 ;
        RECT 242.4375 42.1425 242.7075 42.3675 ;
			LAYER M3 ;
        RECT 242.4375 42.1425 242.7075 42.3675 ;
		END
	END D[11]
	PIN D[12]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
        RECT 242.4375 45.6225 242.7075 45.8475 ;
			LAYER M1 ;
        RECT 242.4375 45.6225 242.7075 45.8475 ;
			LAYER M3 ;
        RECT 242.4375 45.6225 242.7075 45.8475 ;
		END
	END D[12]
	PIN D[13]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
        RECT 242.4375 49.1025 242.7075 49.3275 ;
			LAYER M1 ;
        RECT 242.4375 49.1025 242.7075 49.3275 ;
			LAYER M3 ;
        RECT 242.4375 49.1025 242.7075 49.3275 ;
		END
	END D[13]
	PIN D[14]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
        RECT 242.4375 52.5825 242.7075 52.8075 ;
			LAYER M2 ;
        RECT 242.4375 52.5825 242.7075 52.8075 ;
			LAYER M3 ;
        RECT 242.4375 52.5825 242.7075 52.8075 ;
		END
	END D[14]
	PIN D[15]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
        RECT 242.4375 56.0625 242.7075 56.2875 ;
			LAYER M2 ;
        RECT 242.4375 56.0625 242.7075 56.2875 ;
			LAYER M1 ;
        RECT 242.4375 56.0625 242.7075 56.2875 ;
		END
	END D[15]
	PIN D[16]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
        RECT 242.4375 87.2925 242.7075 87.5175 ;
			LAYER M2 ;
        RECT 242.4375 87.2925 242.7075 87.5175 ;
			LAYER M1 ;
        RECT 242.4375 87.2925 242.7075 87.5175 ;
		END
	END D[16]
	PIN D[17]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
        RECT 242.4375 90.7725 242.7075 90.9975 ;
			LAYER M3 ;
        RECT 242.4375 90.7725 242.7075 90.9975 ;
			LAYER M1 ;
        RECT 242.4375 90.7725 242.7075 90.9975 ;
		END
	END D[17]
	PIN D[18]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
        RECT 242.4375 94.2525 242.7075 94.4775 ;
			LAYER M1 ;
        RECT 242.4375 94.2525 242.7075 94.4775 ;
			LAYER M3 ;
        RECT 242.4375 94.2525 242.7075 94.4775 ;
		END
	END D[18]
	PIN D[19]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
        RECT 242.4375 97.7325 242.7075 97.9575 ;
			LAYER M3 ;
        RECT 242.4375 97.7325 242.7075 97.9575 ;
			LAYER M2 ;
        RECT 242.4375 97.7325 242.7075 97.9575 ;
		END
	END D[19]
	PIN D[1]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
        RECT 242.4375 7.3425 242.7075 7.5675 ;
			LAYER M2 ;
        RECT 242.4375 7.3425 242.7075 7.5675 ;
			LAYER M1 ;
        RECT 242.4375 7.3425 242.7075 7.5675 ;
		END
	END D[1]
	PIN D[20]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
        RECT 242.4375 101.2125 242.7075 101.4375 ;
			LAYER M3 ;
        RECT 242.4375 101.2125 242.7075 101.4375 ;
			LAYER M1 ;
        RECT 242.4375 101.2125 242.7075 101.4375 ;
		END
	END D[20]
	PIN D[21]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
        RECT 242.4375 104.6925 242.7075 104.9175 ;
			LAYER M1 ;
        RECT 242.4375 104.6925 242.7075 104.9175 ;
			LAYER M3 ;
        RECT 242.4375 104.6925 242.7075 104.9175 ;
		END
	END D[21]
	PIN D[22]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
        RECT 242.4375 108.1725 242.7075 108.3975 ;
			LAYER M3 ;
        RECT 242.4375 108.1725 242.7075 108.3975 ;
			LAYER M2 ;
        RECT 242.4375 108.1725 242.7075 108.3975 ;
		END
	END D[22]
	PIN D[23]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
        RECT 242.4375 111.6525 242.7075 111.8775 ;
			LAYER M2 ;
        RECT 242.4375 111.6525 242.7075 111.8775 ;
			LAYER M3 ;
        RECT 242.4375 111.6525 242.7075 111.8775 ;
		END
	END D[23]
	PIN D[24]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
        RECT 242.4375 115.1325 242.7075 115.3575 ;
			LAYER M3 ;
        RECT 242.4375 115.1325 242.7075 115.3575 ;
			LAYER M2 ;
        RECT 242.4375 115.1325 242.7075 115.3575 ;
		END
	END D[24]
	PIN D[25]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
        RECT 242.4375 118.6125 242.7075 118.8375 ;
			LAYER M1 ;
        RECT 242.4375 118.6125 242.7075 118.8375 ;
			LAYER M2 ;
        RECT 242.4375 118.6125 242.7075 118.8375 ;
		END
	END D[25]
	PIN D[26]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
        RECT 242.4375 122.0925 242.7075 122.3175 ;
			LAYER M2 ;
        RECT 242.4375 122.0925 242.7075 122.3175 ;
			LAYER M1 ;
        RECT 242.4375 122.0925 242.7075 122.3175 ;
		END
	END D[26]
	PIN D[27]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
        RECT 242.4375 125.5725 242.7075 125.7975 ;
			LAYER M2 ;
        RECT 242.4375 125.5725 242.7075 125.7975 ;
			LAYER M3 ;
        RECT 242.4375 125.5725 242.7075 125.7975 ;
		END
	END D[27]
	PIN D[28]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
        RECT 242.4375 129.0525 242.7075 129.2775 ;
			LAYER M1 ;
        RECT 242.4375 129.0525 242.7075 129.2775 ;
			LAYER M3 ;
        RECT 242.4375 129.0525 242.7075 129.2775 ;
		END
	END D[28]
	PIN D[29]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
        RECT 242.4375 132.5325 242.7075 132.7575 ;
			LAYER M1 ;
        RECT 242.4375 132.5325 242.7075 132.7575 ;
			LAYER M3 ;
        RECT 242.4375 132.5325 242.7075 132.7575 ;
		END
	END D[29]
	PIN D[2]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
        RECT 242.4375 10.8225 242.7075 11.0475 ;
			LAYER M2 ;
        RECT 242.4375 10.8225 242.7075 11.0475 ;
			LAYER M1 ;
        RECT 242.4375 10.8225 242.7075 11.0475 ;
		END
	END D[2]
	PIN D[30]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
        RECT 242.4375 136.0125 242.7075 136.2375 ;
			LAYER M2 ;
        RECT 242.4375 136.0125 242.7075 136.2375 ;
			LAYER M3 ;
        RECT 242.4375 136.0125 242.7075 136.2375 ;
		END
	END D[30]
	PIN D[31]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
        RECT 242.4375 139.4925 242.7075 139.7175 ;
			LAYER M2 ;
        RECT 242.4375 139.4925 242.7075 139.7175 ;
			LAYER M1 ;
        RECT 242.4375 139.4925 242.7075 139.7175 ;
		END
	END D[31]
	PIN D[3]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
        RECT 242.4375 14.3025 242.7075 14.5275 ;
			LAYER M2 ;
        RECT 242.4375 14.3025 242.7075 14.5275 ;
			LAYER M3 ;
        RECT 242.4375 14.3025 242.7075 14.5275 ;
		END
	END D[3]
	PIN D[4]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
        RECT 242.4375 17.7825 242.7075 18.0075 ;
			LAYER M3 ;
        RECT 242.4375 17.7825 242.7075 18.0075 ;
			LAYER M2 ;
        RECT 242.4375 17.7825 242.7075 18.0075 ;
		END
	END D[4]
	PIN D[5]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
        RECT 242.4375 21.2625 242.7075 21.4875 ;
			LAYER M3 ;
        RECT 242.4375 21.2625 242.7075 21.4875 ;
			LAYER M1 ;
        RECT 242.4375 21.2625 242.7075 21.4875 ;
		END
	END D[5]
	PIN D[6]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
        RECT 242.4375 24.7425 242.7075 24.9675 ;
			LAYER M3 ;
        RECT 242.4375 24.7425 242.7075 24.9675 ;
			LAYER M1 ;
        RECT 242.4375 24.7425 242.7075 24.9675 ;
		END
	END D[6]
	PIN D[7]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
        RECT 242.4375 28.2225 242.7075 28.4475 ;
			LAYER M1 ;
        RECT 242.4375 28.2225 242.7075 28.4475 ;
			LAYER M2 ;
        RECT 242.4375 28.2225 242.7075 28.4475 ;
		END
	END D[7]
	PIN D[8]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
        RECT 242.4375 31.7025 242.7075 31.9275 ;
			LAYER M1 ;
        RECT 242.4375 31.7025 242.7075 31.9275 ;
			LAYER M3 ;
        RECT 242.4375 31.7025 242.7075 31.9275 ;
		END
	END D[8]
	PIN D[9]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
        RECT 242.4375 35.1825 242.7075 35.4075 ;
			LAYER M1 ;
        RECT 242.4375 35.1825 242.7075 35.4075 ;
			LAYER M3 ;
        RECT 242.4375 35.1825 242.7075 35.4075 ;
		END
	END D[9]
	PIN Q[0]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
        RECT 242.4375 2.8950 242.7075 3.1200 ;
			LAYER M3 ;
        RECT 242.4375 2.8950 242.7075 3.1200 ;
			LAYER M2 ;
        RECT 242.4375 2.8950 242.7075 3.1200 ;
		END
	END Q[0]
	PIN Q[10]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
        RECT 242.4375 37.6950 242.7075 37.9200 ;
			LAYER M3 ;
        RECT 242.4375 37.6950 242.7075 37.9200 ;
			LAYER M2 ;
        RECT 242.4375 37.6950 242.7075 37.9200 ;
		END
	END Q[10]
	PIN Q[11]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
        RECT 242.4375 41.1750 242.7075 41.4000 ;
			LAYER M1 ;
        RECT 242.4375 41.1750 242.7075 41.4000 ;
			LAYER M3 ;
        RECT 242.4375 41.1750 242.7075 41.4000 ;
		END
	END Q[11]
	PIN Q[12]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
        RECT 242.4375 44.6550 242.7075 44.8800 ;
			LAYER M1 ;
        RECT 242.4375 44.6550 242.7075 44.8800 ;
			LAYER M2 ;
        RECT 242.4375 44.6550 242.7075 44.8800 ;
		END
	END Q[12]
	PIN Q[13]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
        RECT 242.4375 48.1350 242.7075 48.3600 ;
			LAYER M1 ;
        RECT 242.4375 48.1350 242.7075 48.3600 ;
			LAYER M3 ;
        RECT 242.4375 48.1350 242.7075 48.3600 ;
		END
	END Q[13]
	PIN Q[14]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
        RECT 242.4375 51.6150 242.7075 51.8400 ;
			LAYER M2 ;
        RECT 242.4375 51.6150 242.7075 51.8400 ;
			LAYER M3 ;
        RECT 242.4375 51.6150 242.7075 51.8400 ;
		END
	END Q[14]
	PIN Q[15]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
        RECT 242.4375 55.0950 242.7075 55.3200 ;
			LAYER M1 ;
        RECT 242.4375 55.0950 242.7075 55.3200 ;
			LAYER M3 ;
        RECT 242.4375 55.0950 242.7075 55.3200 ;
		END
	END Q[15]
	PIN Q[16]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
        RECT 242.4375 86.3250 242.7075 86.5500 ;
			LAYER M3 ;
        RECT 242.4375 86.3250 242.7075 86.5500 ;
			LAYER M1 ;
        RECT 242.4375 86.3250 242.7075 86.5500 ;
		END
	END Q[16]
	PIN Q[17]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
        RECT 242.4375 89.8050 242.7075 90.0300 ;
			LAYER M1 ;
        RECT 242.4375 89.8050 242.7075 90.0300 ;
			LAYER M2 ;
        RECT 242.4375 89.8050 242.7075 90.0300 ;
		END
	END Q[17]
	PIN Q[18]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
        RECT 242.4375 93.2850 242.7075 93.5100 ;
			LAYER M1 ;
        RECT 242.4375 93.2850 242.7075 93.5100 ;
			LAYER M3 ;
        RECT 242.4375 93.2850 242.7075 93.5100 ;
		END
	END Q[18]
	PIN Q[19]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
        RECT 242.4375 96.7650 242.7075 96.9900 ;
			LAYER M2 ;
        RECT 242.4375 96.7650 242.7075 96.9900 ;
			LAYER M1 ;
        RECT 242.4375 96.7650 242.7075 96.9900 ;
		END
	END Q[19]
	PIN Q[1]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
        RECT 242.4375 6.3750 242.7075 6.6000 ;
			LAYER M1 ;
        RECT 242.4375 6.3750 242.7075 6.6000 ;
			LAYER M3 ;
        RECT 242.4375 6.3750 242.7075 6.6000 ;
		END
	END Q[1]
	PIN Q[20]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
        RECT 242.4375 100.2450 242.7075 100.4700 ;
			LAYER M3 ;
        RECT 242.4375 100.2450 242.7075 100.4700 ;
			LAYER M1 ;
        RECT 242.4375 100.2450 242.7075 100.4700 ;
		END
	END Q[20]
	PIN Q[21]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
        RECT 242.4375 103.7250 242.7075 103.9500 ;
			LAYER M3 ;
        RECT 242.4375 103.7250 242.7075 103.9500 ;
			LAYER M2 ;
        RECT 242.4375 103.7250 242.7075 103.9500 ;
		END
	END Q[21]
	PIN Q[22]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
        RECT 242.4375 107.2050 242.7075 107.4300 ;
			LAYER M2 ;
        RECT 242.4375 107.2050 242.7075 107.4300 ;
			LAYER M1 ;
        RECT 242.4375 107.2050 242.7075 107.4300 ;
		END
	END Q[22]
	PIN Q[23]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
        RECT 242.4375 110.6850 242.7075 110.9100 ;
			LAYER M3 ;
        RECT 242.4375 110.6850 242.7075 110.9100 ;
			LAYER M1 ;
        RECT 242.4375 110.6850 242.7075 110.9100 ;
		END
	END Q[23]
	PIN Q[24]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
        RECT 242.4375 114.1650 242.7075 114.3900 ;
			LAYER M3 ;
        RECT 242.4375 114.1650 242.7075 114.3900 ;
			LAYER M2 ;
        RECT 242.4375 114.1650 242.7075 114.3900 ;
		END
	END Q[24]
	PIN Q[25]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
        RECT 242.4375 117.6450 242.7075 117.8700 ;
			LAYER M3 ;
        RECT 242.4375 117.6450 242.7075 117.8700 ;
			LAYER M1 ;
        RECT 242.4375 117.6450 242.7075 117.8700 ;
		END
	END Q[25]
	PIN Q[26]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
        RECT 242.4375 121.1250 242.7075 121.3500 ;
			LAYER M1 ;
        RECT 242.4375 121.1250 242.7075 121.3500 ;
			LAYER M2 ;
        RECT 242.4375 121.1250 242.7075 121.3500 ;
		END
	END Q[26]
	PIN Q[27]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
        RECT 242.4375 124.6050 242.7075 124.8300 ;
			LAYER M3 ;
        RECT 242.4375 124.6050 242.7075 124.8300 ;
			LAYER M1 ;
        RECT 242.4375 124.6050 242.7075 124.8300 ;
		END
	END Q[27]
	PIN Q[28]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
        RECT 242.4375 128.0850 242.7075 128.3100 ;
			LAYER M1 ;
        RECT 242.4375 128.0850 242.7075 128.3100 ;
			LAYER M2 ;
        RECT 242.4375 128.0850 242.7075 128.3100 ;
		END
	END Q[28]
	PIN Q[29]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
        RECT 242.4375 131.5650 242.7075 131.7900 ;
			LAYER M1 ;
        RECT 242.4375 131.5650 242.7075 131.7900 ;
			LAYER M3 ;
        RECT 242.4375 131.5650 242.7075 131.7900 ;
		END
	END Q[29]
	PIN Q[2]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
        RECT 242.4375 9.8550 242.7075 10.0800 ;
			LAYER M1 ;
        RECT 242.4375 9.8550 242.7075 10.0800 ;
			LAYER M2 ;
        RECT 242.4375 9.8550 242.7075 10.0800 ;
		END
	END Q[2]
	PIN Q[30]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
        RECT 242.4375 135.0450 242.7075 135.2700 ;
			LAYER M1 ;
        RECT 242.4375 135.0450 242.7075 135.2700 ;
			LAYER M3 ;
        RECT 242.4375 135.0450 242.7075 135.2700 ;
		END
	END Q[30]
	PIN Q[31]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
        RECT 242.4375 138.5250 242.7075 138.7500 ;
			LAYER M1 ;
        RECT 242.4375 138.5250 242.7075 138.7500 ;
			LAYER M3 ;
        RECT 242.4375 138.5250 242.7075 138.7500 ;
		END
	END Q[31]
	PIN Q[3]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
        RECT 242.4375 13.3350 242.7075 13.5600 ;
			LAYER M1 ;
        RECT 242.4375 13.3350 242.7075 13.5600 ;
			LAYER M3 ;
        RECT 242.4375 13.3350 242.7075 13.5600 ;
		END
	END Q[3]
	PIN Q[4]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
        RECT 242.4375 16.8150 242.7075 17.0400 ;
			LAYER M2 ;
        RECT 242.4375 16.8150 242.7075 17.0400 ;
			LAYER M3 ;
        RECT 242.4375 16.8150 242.7075 17.0400 ;
		END
	END Q[4]
	PIN Q[5]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
        RECT 242.4375 20.2950 242.7075 20.5200 ;
			LAYER M3 ;
        RECT 242.4375 20.2950 242.7075 20.5200 ;
			LAYER M2 ;
        RECT 242.4375 20.2950 242.7075 20.5200 ;
		END
	END Q[5]
	PIN Q[6]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
        RECT 242.4375 23.7750 242.7075 24.0000 ;
			LAYER M1 ;
        RECT 242.4375 23.7750 242.7075 24.0000 ;
			LAYER M3 ;
        RECT 242.4375 23.7750 242.7075 24.0000 ;
		END
	END Q[6]
	PIN Q[7]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
        RECT 242.4375 27.2550 242.7075 27.4800 ;
			LAYER M2 ;
        RECT 242.4375 27.2550 242.7075 27.4800 ;
			LAYER M1 ;
        RECT 242.4375 27.2550 242.7075 27.4800 ;
		END
	END Q[7]
	PIN Q[8]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
        RECT 242.4375 30.7350 242.7075 30.9600 ;
			LAYER M2 ;
        RECT 242.4375 30.7350 242.7075 30.9600 ;
			LAYER M3 ;
        RECT 242.4375 30.7350 242.7075 30.9600 ;
		END
	END Q[8]
	PIN Q[9]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
        RECT 242.4375 34.2150 242.7075 34.4400 ;
			LAYER M3 ;
        RECT 242.4375 34.2150 242.7075 34.4400 ;
			LAYER M2 ;
        RECT 242.4375 34.2150 242.7075 34.4400 ;
		END
	END Q[9]
	PIN RTSEL[0]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
        RECT 242.4375 82.8375 242.7075 83.0625 ;
			LAYER M2 ;
        RECT 242.4375 82.8375 242.7075 83.0625 ;
			LAYER M3 ;
        RECT 242.4375 82.8375 242.7075 83.0625 ;
		END
	END RTSEL[0]
	PIN RTSEL[1]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
        RECT 242.4375 83.3325 242.7075 83.5575 ;
			LAYER M2 ;
        RECT 242.4375 83.3325 242.7075 83.5575 ;
			LAYER M3 ;
        RECT 242.4375 83.3325 242.7075 83.5575 ;
		END
	END RTSEL[1]
	PIN SD
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
        RECT 242.4375 77.0325 242.7075 77.2575 ;
			LAYER M1 ;
        RECT 242.4375 77.0325 242.7075 77.2575 ;
			LAYER M3 ;
        RECT 242.4375 77.0325 242.7075 77.2575 ;
		END
	END SD
	PIN SLP
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
        RECT 242.4375 76.4475 242.7075 76.6725 ;
			LAYER M3 ;
        RECT 242.4375 76.4475 242.7075 76.6725 ;
			LAYER M1 ;
        RECT 242.4375 76.4475 242.7075 76.6725 ;
		END
	END SLP
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M4 ;
        RECT 0.0000 4.2225 242.1300 4.6575 ;
			LAYER M4 ;
        RECT 0.0000 7.7025 242.1300 8.1375 ;
			LAYER M4 ;
        RECT 0.0000 11.1825 242.1300 11.6175 ;
			LAYER M4 ;
        RECT 0.0000 14.6625 242.1300 15.0975 ;
			LAYER M4 ;
        RECT 0.0000 18.1425 242.1300 18.5775 ;
			LAYER M4 ;
        RECT 0.0000 21.6225 242.1300 22.0575 ;
			LAYER M4 ;
        RECT 0.0000 25.1025 242.1300 25.5375 ;
			LAYER M4 ;
        RECT 0.0000 28.5825 242.1300 29.0175 ;
			LAYER M4 ;
        RECT 0.0000 32.0625 242.1300 32.4975 ;
			LAYER M4 ;
        RECT 0.0000 35.5425 242.1300 35.9775 ;
			LAYER M4 ;
        RECT 0.0000 39.0225 242.1300 39.4575 ;
			LAYER M4 ;
        RECT 0.0000 42.5025 242.1300 42.9375 ;
			LAYER M4 ;
        RECT 0.0000 45.9825 242.1300 46.4175 ;
			LAYER M4 ;
        RECT 0.0000 49.4625 242.1300 49.8975 ;
			LAYER M4 ;
        RECT 0.0000 52.9425 242.1300 53.3775 ;
			LAYER M4 ;
        RECT 0.0000 56.4225 242.1300 56.8575 ;
			LAYER M4 ;
        RECT 0.0000 59.6325 242.2050 60.2625 ;
			LAYER M4 ;
        RECT 0.0000 64.5375 242.2050 65.1675 ;
			LAYER M4 ;
        RECT 0.0000 75.6375 242.2050 76.2675 ;
			LAYER M4 ;
        RECT 0.0000 80.9250 242.2050 81.5550 ;
			LAYER M4 ;
        RECT 0.0000 87.6525 242.1300 88.0875 ;
			LAYER M4 ;
        RECT 0.0000 91.1325 242.1300 91.5675 ;
			LAYER M4 ;
        RECT 0.0000 94.6125 242.1300 95.0475 ;
			LAYER M4 ;
        RECT 0.0000 98.0925 242.1300 98.5275 ;
			LAYER M4 ;
        RECT 0.0000 101.5725 242.1300 102.0075 ;
			LAYER M4 ;
        RECT 0.0000 105.0525 242.1300 105.4875 ;
			LAYER M4 ;
        RECT 0.0000 108.5325 242.1300 108.9675 ;
			LAYER M4 ;
        RECT 0.0000 112.0125 242.1300 112.4475 ;
			LAYER M4 ;
        RECT 0.0000 115.4925 242.1300 115.9275 ;
			LAYER M4 ;
        RECT 0.0000 118.9725 242.1300 119.4075 ;
			LAYER M4 ;
        RECT 0.0000 122.4525 242.1300 122.8875 ;
			LAYER M4 ;
        RECT 0.0000 125.9325 242.1300 126.3675 ;
			LAYER M4 ;
        RECT 0.0000 129.4125 242.1300 129.8475 ;
			LAYER M4 ;
        RECT 0.0000 132.8925 242.1300 133.3275 ;
			LAYER M4 ;
        RECT 0.0000 136.3725 242.1300 136.8075 ;
			LAYER M4 ;
        RECT 0.0000 139.8525 242.1300 140.2875 ;
		END
	END VDD
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M4 ;
        RECT 0.0000 1.3275 242.1300 1.7625 ;
			LAYER M4 ;
        RECT 0.0000 4.8075 242.1300 5.2425 ;
			LAYER M4 ;
        RECT 0.0000 8.2875 242.1300 8.7225 ;
			LAYER M4 ;
        RECT 0.0000 11.7675 242.1300 12.2025 ;
			LAYER M4 ;
        RECT 0.0000 15.2475 242.1300 15.6825 ;
			LAYER M4 ;
        RECT 0.0000 18.7275 242.1300 19.1625 ;
			LAYER M4 ;
        RECT 0.0000 22.2075 242.1300 22.6425 ;
			LAYER M4 ;
        RECT 0.0000 25.6875 242.1300 26.1225 ;
			LAYER M4 ;
        RECT 0.0000 29.1675 242.1300 29.6025 ;
			LAYER M4 ;
        RECT 0.0000 32.6475 242.1300 33.0825 ;
			LAYER M4 ;
        RECT 0.0000 36.1275 242.1300 36.5625 ;
			LAYER M4 ;
        RECT 0.0000 39.6075 242.1300 40.0425 ;
			LAYER M4 ;
        RECT 0.0000 43.0875 242.1300 43.5225 ;
			LAYER M4 ;
        RECT 0.0000 46.5675 242.1300 47.0025 ;
			LAYER M4 ;
        RECT 0.0000 50.0475 242.1300 50.4825 ;
			LAYER M4 ;
        RECT 0.0000 53.5275 242.1300 53.9625 ;
			LAYER M4 ;
        RECT 0.0000 62.0025 242.2050 62.6325 ;
			LAYER M4 ;
        RECT 0.0000 68.1750 242.2050 68.8050 ;
			LAYER M4 ;
        RECT 0.0000 72.6075 242.2050 73.2375 ;
			LAYER M4 ;
        RECT 0.0000 77.6925 242.2050 78.3225 ;
			LAYER M4 ;
        RECT 0.0000 84.7575 242.1300 85.1925 ;
			LAYER M4 ;
        RECT 0.0000 88.2375 242.1300 88.6725 ;
			LAYER M4 ;
        RECT 0.0000 91.7175 242.1300 92.1525 ;
			LAYER M4 ;
        RECT 0.0000 95.1975 242.1300 95.6325 ;
			LAYER M4 ;
        RECT 0.0000 98.6775 242.1300 99.1125 ;
			LAYER M4 ;
        RECT 0.0000 102.1575 242.1300 102.5925 ;
			LAYER M4 ;
        RECT 0.0000 105.6375 242.1300 106.0725 ;
			LAYER M4 ;
        RECT 0.0000 109.1175 242.1300 109.5525 ;
			LAYER M4 ;
        RECT 0.0000 112.5975 242.1300 113.0325 ;
			LAYER M4 ;
        RECT 0.0000 116.0775 242.1300 116.5125 ;
			LAYER M4 ;
        RECT 0.0000 119.5575 242.1300 119.9925 ;
			LAYER M4 ;
        RECT 0.0000 123.0375 242.1300 123.4725 ;
			LAYER M4 ;
        RECT 0.0000 126.5175 242.1300 126.9525 ;
			LAYER M4 ;
        RECT 0.0000 129.9975 242.1300 130.4325 ;
			LAYER M4 ;
        RECT 0.0000 133.4775 242.1300 133.9125 ;
			LAYER M4 ;
        RECT 0.0000 136.9575 242.1300 137.3925 ;
		END
	END VSS
	PIN WEB
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
        RECT 242.4375 64.5900 242.7075 64.8150 ;
			LAYER M1 ;
        RECT 242.4375 64.5900 242.7075 64.8150 ;
			LAYER M3 ;
        RECT 242.4375 64.5900 242.7075 64.8150 ;
		END
	END WEB
	PIN WEBM
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
        RECT 242.4375 65.2800 242.7075 65.5050 ;
			LAYER M2 ;
        RECT 242.4375 65.2800 242.7075 65.5050 ;
			LAYER M1 ;
        RECT 242.4375 65.2800 242.7075 65.5050 ;
		END
	END WEBM
	PIN WTSEL[0]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
        RECT 242.4375 81.7050 242.7075 81.9300 ;
			LAYER M1 ;
        RECT 242.4375 81.7050 242.7075 81.9300 ;
			LAYER M2 ;
        RECT 242.4375 81.7050 242.7075 81.9300 ;
		END
	END WTSEL[0]
	PIN WTSEL[1]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
        RECT 242.4375 83.8275 242.7075 84.0525 ;
			LAYER M2 ;
        RECT 242.4375 83.8275 242.7075 84.0525 ;
			LAYER M3 ;
        RECT 242.4375 83.8275 242.7075 84.0525 ;
		END
	END WTSEL[1]
	OBS
		LAYER M2 ;
        RECT 242.4375 11.6625 242.7075 11.7225 ;
		LAYER M1 ;
        RECT 242.4375 18.5925 242.7075 18.7125 ;
		LAYER M3 ;
        RECT 242.4375 18.1275 242.7075 18.1575 ;
		LAYER M3 ;
        RECT 242.4375 41.5200 242.7075 42.0225 ;
		LAYER M2 ;
        RECT 242.4375 58.4400 242.7075 58.4700 ;
		LAYER M1 ;
        RECT 242.4375 58.4100 242.7075 58.5000 ;
		LAYER M3 ;
        RECT 242.4375 58.9350 242.7075 58.9650 ;
		LAYER M1 ;
        RECT 242.4375 49.9125 242.7075 50.0325 ;
		LAYER VIA3 ;
        RECT 242.4375 58.9350 242.7075 58.9650 ;
		LAYER VIA3 ;
        RECT 242.4375 52.9275 242.7075 52.9575 ;
		LAYER M3 ;
        RECT 242.4375 53.9475 242.7075 53.9775 ;
		LAYER VIA3 ;
        RECT 242.4375 49.9425 242.7075 50.0025 ;
		LAYER M2 ;
        RECT 242.4375 49.9425 242.7075 50.0025 ;
		LAYER M2 ;
        RECT 242.4375 52.9275 242.7075 52.9575 ;
		LAYER VIA3 ;
        RECT 242.4375 58.4400 242.7075 58.4700 ;
		LAYER M3 ;
        RECT 242.4375 56.9025 242.7075 57.9750 ;
		LAYER VIA3 ;
        RECT 242.4375 56.9025 242.7075 57.9750 ;
		LAYER M3 ;
        RECT 242.4375 55.4400 242.7075 55.9425 ;
		LAYER M2 ;
        RECT 242.4375 56.9025 242.7075 57.9750 ;
		LAYER M3 ;
        RECT 242.4375 19.6425 242.7075 20.1750 ;
		LAYER M2 ;
        RECT 242.4375 19.6425 242.7075 20.1750 ;
		LAYER M2 ;
        RECT 242.4375 18.6225 242.7075 18.6825 ;
		LAYER M3 ;
        RECT 242.4375 18.6225 242.7075 18.6825 ;
		LAYER VIA3 ;
        RECT 242.4375 18.6225 242.7075 18.6825 ;
		LAYER VIA3 ;
        RECT 242.4375 34.5600 242.7075 35.0625 ;
		LAYER M3 ;
        RECT 242.4375 25.5825 242.7075 25.6425 ;
		LAYER M1 ;
        RECT 242.4375 25.5525 242.7075 25.6725 ;
		LAYER VIA3 ;
        RECT 242.4375 26.6025 242.7075 27.1350 ;
		LAYER M2 ;
        RECT 242.4375 26.6025 242.7075 27.1350 ;
		LAYER M1 ;
        RECT 242.4375 29.0325 242.7075 29.1525 ;
		LAYER M3 ;
        RECT 242.4375 30.0825 242.7075 30.6150 ;
		LAYER M2 ;
        RECT 242.4375 29.5875 242.7075 29.6175 ;
		LAYER M1 ;
        RECT 242.4375 29.5575 242.7075 29.6475 ;
		LAYER M2 ;
        RECT 242.4375 28.5675 242.7075 28.5975 ;
		LAYER M3 ;
        RECT 242.4375 28.5675 242.7075 28.5975 ;
		LAYER M1 ;
        RECT 242.4375 28.5375 242.7075 28.6275 ;
		LAYER VIA3 ;
        RECT 242.4375 27.6000 242.7075 28.1025 ;
		LAYER VIA3 ;
        RECT 242.4375 28.5675 242.7075 28.5975 ;
		LAYER VIA3 ;
        RECT 242.4375 40.0275 242.7075 40.0575 ;
		LAYER M2 ;
        RECT 242.4375 39.5025 242.7075 39.5625 ;
		LAYER VIA3 ;
        RECT 242.4375 39.5025 242.7075 39.5625 ;
		LAYER M3 ;
        RECT 242.4375 39.5025 242.7075 39.5625 ;
		LAYER VIA3 ;
        RECT 242.4375 39.0075 242.7075 39.0375 ;
		LAYER M1 ;
        RECT 242.4375 38.9775 242.7075 39.0675 ;
		LAYER VIA3 ;
        RECT 242.4375 38.0400 242.7075 38.5425 ;
		LAYER M3 ;
        RECT 242.4375 38.0400 242.7075 38.5425 ;
		LAYER M2 ;
        RECT 242.4375 37.0425 242.7075 37.5750 ;
		LAYER M3 ;
        RECT 242.4375 37.0425 242.7075 37.5750 ;
		LAYER VIA3 ;
        RECT 242.4375 37.0425 242.7075 37.5750 ;
		LAYER VIA3 ;
        RECT 242.4375 36.5475 242.7075 36.5775 ;
		LAYER M1 ;
        RECT 242.4375 37.0125 242.7075 37.6050 ;
		LAYER M1 ;
        RECT 242.4375 36.5175 242.7075 36.6075 ;
		LAYER M1 ;
        RECT 242.4375 35.4975 242.7075 35.5875 ;
		LAYER M2 ;
        RECT 242.4375 36.5475 242.7075 36.5775 ;
		LAYER M3 ;
        RECT 242.4375 36.5475 242.7075 36.5775 ;
		LAYER M1 ;
        RECT 242.4375 35.9925 242.7075 36.1125 ;
		LAYER M2 ;
        RECT 242.4375 40.0275 242.7075 40.0575 ;
		LAYER M3 ;
        RECT 242.4375 40.0275 242.7075 40.0575 ;
		LAYER M1 ;
        RECT 242.4375 39.4725 242.7075 39.5925 ;
		LAYER M2 ;
        RECT 242.4375 39.0075 242.7075 39.0375 ;
		LAYER M3 ;
        RECT 242.4375 39.0075 242.7075 39.0375 ;
		LAYER M2 ;
        RECT 242.4375 38.0400 242.7075 38.5425 ;
		LAYER M2 ;
        RECT 242.4375 34.5600 242.7075 35.0625 ;
		LAYER M2 ;
        RECT 242.4375 32.5425 242.7075 32.6025 ;
		LAYER VIA3 ;
        RECT 242.4375 33.0675 242.7075 33.0975 ;
		LAYER M1 ;
        RECT 242.4375 33.0375 242.7075 33.1275 ;
		LAYER M1 ;
        RECT 242.4375 32.5125 242.7075 32.6325 ;
		LAYER M2 ;
        RECT 242.4375 32.0475 242.7075 32.0775 ;
		LAYER VIA3 ;
        RECT 242.4375 32.0475 242.7075 32.0775 ;
		LAYER M1 ;
        RECT 242.4375 32.0175 242.7075 32.1075 ;
		LAYER VIA3 ;
        RECT 242.4375 31.0800 242.7075 31.5825 ;
		LAYER M2 ;
        RECT 242.4375 31.0800 242.7075 31.5825 ;
		LAYER M1 ;
        RECT 242.4375 31.0500 242.7075 31.6125 ;
		LAYER M3 ;
        RECT 242.4375 32.5425 242.7075 32.6025 ;
		LAYER VIA3 ;
        RECT 242.4375 30.0825 242.7075 30.6150 ;
		LAYER M2 ;
        RECT 242.4375 30.0825 242.7075 30.6150 ;
		LAYER M1 ;
        RECT 242.4375 41.4900 242.7075 42.0525 ;
		LAYER M2 ;
        RECT 242.4375 42.9825 242.7075 43.0425 ;
		LAYER VIA3 ;
        RECT 242.4375 44.0025 242.7075 44.5350 ;
		LAYER M2 ;
        RECT 242.4375 45.9675 242.7075 45.9975 ;
		LAYER M3 ;
        RECT 242.4375 43.5075 242.7075 43.5375 ;
		LAYER M1 ;
        RECT 242.4375 42.4575 242.7075 42.5475 ;
		LAYER M2 ;
        RECT 242.4375 40.5225 242.7075 41.0550 ;
		LAYER M3 ;
        RECT 242.4375 40.5225 242.7075 41.0550 ;
		LAYER M2 ;
        RECT 242.4375 47.4825 242.7075 48.0150 ;
		LAYER M2 ;
        RECT 242.4375 41.5200 242.7075 42.0225 ;
		LAYER M3 ;
        RECT 242.4375 47.4825 242.7075 48.0150 ;
		LAYER M3 ;
        RECT 242.4375 49.4475 242.7075 49.4775 ;
		LAYER M1 ;
        RECT 242.4375 49.4175 242.7075 49.5075 ;
		LAYER VIA3 ;
        RECT 242.4375 48.4800 242.7075 48.9825 ;
		LAYER M3 ;
        RECT 242.4375 35.5275 242.7075 35.5575 ;
		LAYER M1 ;
        RECT 242.4375 39.9975 242.7075 40.0875 ;
		LAYER M1 ;
        RECT 242.4375 38.0100 242.7075 38.5725 ;
		LAYER M1 ;
        RECT 242.4375 40.4925 242.7075 41.0850 ;
		LAYER M3 ;
        RECT 242.4375 46.4625 242.7075 46.5225 ;
		LAYER M2 ;
        RECT 242.4375 46.9875 242.7075 47.0175 ;
		LAYER M3 ;
        RECT 242.4375 46.9875 242.7075 47.0175 ;
		LAYER VIA3 ;
        RECT 242.4375 40.5225 242.7075 41.0550 ;
		LAYER M3 ;
        RECT 242.4375 72.2550 242.7075 72.4800 ;
		LAYER M1 ;
        RECT 242.4375 72.2250 242.7075 72.5100 ;
		LAYER M2 ;
        RECT 242.4375 72.9450 242.7075 72.9750 ;
		LAYER VIA3 ;
        RECT 242.4375 72.9450 242.7075 72.9750 ;
		LAYER M2 ;
        RECT 242.4375 74.1300 242.7075 74.6250 ;
		LAYER M3 ;
        RECT 242.4375 74.1300 242.7075 74.6250 ;
		LAYER VIA3 ;
        RECT 242.4375 74.1300 242.7075 74.6250 ;
		LAYER M1 ;
        RECT 242.4375 70.5750 242.7075 70.8600 ;
		LAYER M1 ;
        RECT 242.4375 70.0800 242.7075 70.1700 ;
		LAYER M1 ;
        RECT 242.4375 71.2650 242.7075 71.8200 ;
		LAYER M2 ;
        RECT 242.4375 73.4400 242.7075 73.6650 ;
		LAYER M1 ;
        RECT 242.4375 68.4300 242.7075 68.9850 ;
		LAYER VIA3 ;
        RECT 242.4375 69.4200 242.7075 69.6450 ;
		LAYER M1 ;
        RECT 242.4375 69.3900 242.7075 69.6750 ;
		LAYER M1 ;
        RECT 242.4375 67.7400 242.7075 68.0250 ;
		LAYER VIA3 ;
        RECT 242.4375 70.6050 242.7075 70.8300 ;
		LAYER M1 ;
        RECT 242.4375 73.4100 242.7075 73.6950 ;
		LAYER M3 ;
        RECT 242.4375 73.4400 242.7075 73.6650 ;
		LAYER M2 ;
        RECT 242.4375 70.6050 242.7075 70.8300 ;
		LAYER M3 ;
        RECT 242.4375 70.6050 242.7075 70.8300 ;
		LAYER VIA3 ;
        RECT 242.4375 72.2550 242.7075 72.4800 ;
		LAYER VIA3 ;
        RECT 242.4375 71.2950 242.7075 71.7900 ;
		LAYER M3 ;
        RECT 242.4375 71.2950 242.7075 71.7900 ;
		LAYER M2 ;
        RECT 242.4375 124.9500 242.7075 125.4525 ;
		LAYER M2 ;
        RECT 242.4375 122.4375 242.7075 122.4675 ;
		LAYER M3 ;
        RECT 242.4375 122.4375 242.7075 122.4675 ;
		LAYER M1 ;
        RECT 242.4375 123.9225 242.7075 124.5150 ;
		LAYER VIA3 ;
        RECT 242.4375 122.4375 242.7075 122.4675 ;
		LAYER M3 ;
        RECT 242.4375 123.9525 242.7075 124.4850 ;
		LAYER M2 ;
        RECT 242.4375 122.9325 242.7075 122.9925 ;
		LAYER M3 ;
        RECT 242.4375 122.9325 242.7075 122.9925 ;
		LAYER VIA3 ;
        RECT 242.4375 122.9325 242.7075 122.9925 ;
		LAYER M2 ;
        RECT 242.4375 123.9525 242.7075 124.4850 ;
		LAYER M3 ;
        RECT 242.4375 113.0175 242.7075 113.0475 ;
		LAYER VIA3 ;
        RECT 242.4375 113.0175 242.7075 113.0475 ;
		LAYER M2 ;
        RECT 242.4375 113.0175 242.7075 113.0475 ;
		LAYER M2 ;
        RECT 242.4375 112.4925 242.7075 112.5525 ;
		LAYER VIA3 ;
        RECT 242.4375 112.4925 242.7075 112.5525 ;
		LAYER M1 ;
        RECT 242.4375 112.9875 242.7075 113.0775 ;
		LAYER M3 ;
        RECT 242.4375 124.9500 242.7075 125.4525 ;
		LAYER M2 ;
        RECT 242.4375 120.4725 242.7075 121.0050 ;
		LAYER VIA3 ;
        RECT 242.4375 123.9525 242.7075 124.4850 ;
		LAYER M3 ;
        RECT 242.4375 121.4700 242.7075 121.9725 ;
		LAYER VIA3 ;
        RECT 242.4375 121.4700 242.7075 121.9725 ;
		LAYER M1 ;
        RECT 242.4375 121.4400 242.7075 122.0025 ;
		LAYER M1 ;
        RECT 242.4375 122.4075 242.7075 122.4975 ;
		LAYER M3 ;
        RECT 242.4375 119.9775 242.7075 120.0075 ;
		LAYER VIA3 ;
        RECT 242.4375 119.9775 242.7075 120.0075 ;
		LAYER VIA3 ;
        RECT 242.4375 118.9575 242.7075 118.9875 ;
		LAYER M2 ;
        RECT 242.4375 117.9900 242.7075 118.4925 ;
		LAYER M2 ;
        RECT 242.4375 119.9775 242.7075 120.0075 ;
		LAYER VIA3 ;
        RECT 242.4375 124.9500 242.7075 125.4525 ;
		LAYER M3 ;
        RECT 242.4375 112.4925 242.7075 112.5525 ;
		LAYER M1 ;
        RECT 242.4375 119.9475 242.7075 120.0375 ;
		LAYER M1 ;
        RECT 242.4375 120.4425 242.7075 121.0350 ;
		LAYER M1 ;
        RECT 242.4375 112.4625 242.7075 112.5825 ;
		LAYER M1 ;
        RECT 242.4375 111.9675 242.7075 112.0575 ;
		LAYER M2 ;
        RECT 242.4375 116.4975 242.7075 116.5275 ;
		LAYER M3 ;
        RECT 242.4375 116.4975 242.7075 116.5275 ;
		LAYER VIA3 ;
        RECT 242.4375 115.9725 242.7075 116.0325 ;
		LAYER VIA3 ;
        RECT 242.4375 116.4975 242.7075 116.5275 ;
		LAYER M3 ;
        RECT 242.4375 115.9725 242.7075 116.0325 ;
		LAYER M2 ;
        RECT 242.4375 115.9725 242.7075 116.0325 ;
		LAYER M3 ;
        RECT 242.4375 114.5100 242.7075 115.0125 ;
		LAYER M1 ;
        RECT 242.4375 114.4800 242.7075 115.0425 ;
		LAYER M3 ;
        RECT 242.4375 115.4775 242.7075 115.5075 ;
		LAYER VIA3 ;
        RECT 242.4375 115.4775 242.7075 115.5075 ;
		LAYER M3 ;
        RECT 242.4375 113.5125 242.7075 114.0450 ;
		LAYER M1 ;
        RECT 242.4375 117.9600 242.7075 118.5225 ;
		LAYER VIA3 ;
        RECT 242.4375 117.9900 242.7075 118.4925 ;
		LAYER M1 ;
        RECT 242.4375 116.9625 242.7075 117.5550 ;
		LAYER M1 ;
        RECT 242.4375 113.4825 242.7075 114.0750 ;
		LAYER VIA3 ;
        RECT 242.4375 113.5125 242.7075 114.0450 ;
		LAYER M2 ;
        RECT 242.4375 113.5125 242.7075 114.0450 ;
		LAYER M1 ;
        RECT 242.4375 115.9425 242.7075 116.0625 ;
		LAYER M1 ;
        RECT 242.4375 116.4675 242.7075 116.5575 ;
		LAYER M1 ;
        RECT 242.4375 115.4475 242.7075 115.5375 ;
		LAYER VIA3 ;
        RECT 242.4375 116.9925 242.7075 117.5250 ;
		LAYER M3 ;
        RECT 242.4375 116.9925 242.7075 117.5250 ;
		LAYER M2 ;
        RECT 242.4375 116.9925 242.7075 117.5250 ;
		LAYER M2 ;
        RECT 242.4375 114.5100 242.7075 115.0125 ;
		LAYER VIA3 ;
        RECT 242.4375 114.5100 242.7075 115.0125 ;
		LAYER M2 ;
        RECT 242.4375 115.4775 242.7075 115.5075 ;
		LAYER M3 ;
        RECT 242.4375 11.6625 242.7075 11.7225 ;
		LAYER M3 ;
        RECT 242.4375 13.6800 242.7075 14.1825 ;
		LAYER VIA3 ;
        RECT 242.4375 14.6475 242.7075 14.6775 ;
		LAYER M1 ;
        RECT 242.4375 13.6500 242.7075 14.2125 ;
		LAYER VIA3 ;
        RECT 242.4375 11.6625 242.7075 11.7225 ;
		LAYER M1 ;
        RECT 242.4375 12.1575 242.7075 12.2475 ;
		LAYER M2 ;
        RECT 242.4375 12.1875 242.7075 12.2175 ;
		LAYER M3 ;
        RECT 242.4375 12.6825 242.7075 13.2150 ;
		LAYER M1 ;
        RECT 242.4375 12.6525 242.7075 13.2450 ;
		LAYER M2 ;
        RECT 242.4375 13.6800 242.7075 14.1825 ;
		LAYER M2 ;
        RECT 242.4375 12.6825 242.7075 13.2150 ;
		LAYER VIA3 ;
        RECT 242.4375 12.6825 242.7075 13.2150 ;
		LAYER M2 ;
        RECT 242.4375 25.0875 242.7075 25.1175 ;
		LAYER M3 ;
        RECT 242.4375 22.1025 242.7075 22.1625 ;
		LAYER VIA3 ;
        RECT 242.4375 22.1025 242.7075 22.1625 ;
		LAYER M3 ;
        RECT 242.4375 12.1875 242.7075 12.2175 ;
		LAYER VIA3 ;
        RECT 242.4375 12.1875 242.7075 12.2175 ;
		LAYER VIA3 ;
        RECT 242.4375 13.6800 242.7075 14.1825 ;
		LAYER M1 ;
        RECT 242.4375 18.0975 242.7075 18.1875 ;
		LAYER M2 ;
        RECT 242.4375 18.1275 242.7075 18.1575 ;
		LAYER VIA3 ;
        RECT 242.4375 18.1275 242.7075 18.1575 ;
		LAYER M3 ;
        RECT 242.4375 16.1625 242.7075 16.6950 ;
		LAYER VIA3 ;
        RECT 242.4375 16.1625 242.7075 16.6950 ;
		LAYER M1 ;
        RECT 242.4375 16.1325 242.7075 16.7250 ;
		LAYER M2 ;
        RECT 242.4375 16.1625 242.7075 16.6950 ;
		LAYER VIA3 ;
        RECT 242.4375 20.6400 242.7075 21.1425 ;
		LAYER M1 ;
        RECT 242.4375 19.6125 242.7075 20.2050 ;
		LAYER VIA3 ;
        RECT 242.4375 19.1475 242.7075 19.1775 ;
		LAYER M3 ;
        RECT 242.4375 19.1475 242.7075 19.1775 ;
		LAYER M3 ;
        RECT 242.4375 20.6400 242.7075 21.1425 ;
		LAYER M2 ;
        RECT 242.4375 20.6400 242.7075 21.1425 ;
		LAYER M2 ;
        RECT 242.4375 19.1475 242.7075 19.1775 ;
		LAYER M1 ;
        RECT 242.4375 19.1175 242.7075 19.2075 ;
		LAYER M3 ;
        RECT 242.4375 17.1600 242.7075 17.6625 ;
		LAYER VIA3 ;
        RECT 242.4375 17.1600 242.7075 17.6625 ;
		LAYER M2 ;
        RECT 242.4375 17.1600 242.7075 17.6625 ;
		LAYER M1 ;
        RECT 242.4375 17.1300 242.7075 17.6925 ;
		LAYER M1 ;
        RECT 242.4375 34.5300 242.7075 35.0925 ;
		LAYER M3 ;
        RECT 242.4375 34.5600 242.7075 35.0625 ;
		LAYER M1 ;
        RECT 242.4375 30.0525 242.7075 30.6450 ;
		LAYER VIA3 ;
        RECT 242.4375 33.5625 242.7075 34.0950 ;
		LAYER M3 ;
        RECT 242.4375 33.5625 242.7075 34.0950 ;
		LAYER M2 ;
        RECT 242.4375 33.5625 242.7075 34.0950 ;
		LAYER M1 ;
        RECT 242.4375 33.5325 242.7075 34.1250 ;
		LAYER VIA3 ;
        RECT 242.4375 36.0225 242.7075 36.0825 ;
		LAYER M3 ;
        RECT 242.4375 36.0225 242.7075 36.0825 ;
		LAYER M2 ;
        RECT 242.4375 35.5275 242.7075 35.5575 ;
		LAYER VIA3 ;
        RECT 242.4375 35.5275 242.7075 35.5575 ;
		LAYER M2 ;
        RECT 242.4375 36.0225 242.7075 36.0825 ;
		LAYER M2 ;
        RECT 242.4375 33.0675 242.7075 33.0975 ;
		LAYER M3 ;
        RECT 242.4375 33.0675 242.7075 33.0975 ;
		LAYER M3 ;
        RECT 242.4375 32.0475 242.7075 32.0775 ;
		LAYER M3 ;
        RECT 242.4375 31.0800 242.7075 31.5825 ;
		LAYER VIA3 ;
        RECT 242.4375 32.5425 242.7075 32.6025 ;
		LAYER M1 ;
        RECT 242.4375 15.6375 242.7075 15.7275 ;
		LAYER M2 ;
        RECT 242.4375 15.1425 242.7075 15.2025 ;
		LAYER M1 ;
        RECT 242.4375 15.1125 242.7075 15.2325 ;
		LAYER M3 ;
        RECT 242.4375 15.1425 242.7075 15.2025 ;
		LAYER VIA3 ;
        RECT 242.4375 15.1425 242.7075 15.2025 ;
		LAYER M3 ;
        RECT 242.4375 15.6675 242.7075 15.6975 ;
		LAYER M2 ;
        RECT 242.4375 24.1200 242.7075 24.6225 ;
		LAYER VIA3 ;
        RECT 242.4375 24.1200 242.7075 24.6225 ;
		LAYER M1 ;
        RECT 242.4375 25.0575 242.7075 25.1475 ;
		LAYER M1 ;
        RECT 242.4375 26.0775 242.7075 26.1675 ;
		LAYER M3 ;
        RECT 242.4375 24.1200 242.7075 24.6225 ;
		LAYER M1 ;
        RECT 242.4375 27.5700 242.7075 28.1325 ;
		LAYER M2 ;
        RECT 242.4375 29.0625 242.7075 29.1225 ;
		LAYER M3 ;
        RECT 242.4375 29.0625 242.7075 29.1225 ;
		LAYER M3 ;
        RECT 242.4375 29.5875 242.7075 29.6175 ;
		LAYER M2 ;
        RECT 242.4375 27.6000 242.7075 28.1025 ;
		LAYER VIA3 ;
        RECT 242.4375 29.0625 242.7075 29.1225 ;
		LAYER M3 ;
        RECT 242.4375 27.6000 242.7075 28.1025 ;
		LAYER VIA3 ;
        RECT 242.4375 29.5875 242.7075 29.6175 ;
		LAYER M1 ;
        RECT 242.4375 26.5725 242.7075 27.1650 ;
		LAYER M3 ;
        RECT 242.4375 26.6025 242.7075 27.1350 ;
		LAYER M1 ;
        RECT 242.4375 20.6100 242.7075 21.1725 ;
		LAYER M2 ;
        RECT 242.4375 21.6075 242.7075 21.6375 ;
		LAYER M1 ;
        RECT 242.4375 21.5775 242.7075 21.6675 ;
		LAYER VIA3 ;
        RECT 242.4375 19.6425 242.7075 20.1750 ;
		LAYER M3 ;
        RECT 242.4375 21.6075 242.7075 21.6375 ;
		LAYER VIA3 ;
        RECT 242.4375 21.6075 242.7075 21.6375 ;
		LAYER M3 ;
        RECT 242.4375 22.6275 242.7075 22.6575 ;
		LAYER M2 ;
        RECT 242.4375 22.6275 242.7075 22.6575 ;
		LAYER M1 ;
        RECT 242.4375 22.5975 242.7075 22.6875 ;
		LAYER M2 ;
        RECT 242.4375 22.1025 242.7075 22.1625 ;
		LAYER M1 ;
        RECT 242.4375 22.0725 242.7075 22.1925 ;
		LAYER VIA3 ;
        RECT 242.4375 22.6275 242.7075 22.6575 ;
		LAYER VIA3 ;
        RECT 242.4375 23.1225 242.7075 23.6550 ;
		LAYER M3 ;
        RECT 242.4375 23.1225 242.7075 23.6550 ;
		LAYER M1 ;
        RECT 242.4375 24.0900 242.7075 24.6525 ;
		LAYER M2 ;
        RECT 242.4375 23.1225 242.7075 23.6550 ;
		LAYER M1 ;
        RECT 242.4375 23.0925 242.7075 23.6850 ;
		LAYER M3 ;
        RECT 242.4375 25.0875 242.7075 25.1175 ;
		LAYER M2 ;
        RECT 242.4375 25.5825 242.7075 25.6425 ;
		LAYER VIA3 ;
        RECT 242.4375 25.5825 242.7075 25.6425 ;
		LAYER M3 ;
        RECT 242.4375 26.1075 242.7075 26.1375 ;
		LAYER VIA3 ;
        RECT 242.4375 25.0875 242.7075 25.1175 ;
		LAYER M2 ;
        RECT 242.4375 26.1075 242.7075 26.1375 ;
		LAYER VIA3 ;
        RECT 242.4375 26.1075 242.7075 26.1375 ;
		LAYER VIA3 ;
        RECT 242.4375 68.4600 242.7075 68.9550 ;
		LAYER M2 ;
        RECT 242.4375 75.0900 242.7075 75.3150 ;
		LAYER M3 ;
        RECT 242.4375 75.0900 242.7075 75.3150 ;
		LAYER VIA3 ;
        RECT 242.4375 75.0900 242.7075 75.3150 ;
		LAYER VIA3 ;
        RECT 242.4375 73.4400 242.7075 73.6650 ;
		LAYER M2 ;
        RECT 242.4375 71.2950 242.7075 71.7900 ;
		LAYER M3 ;
        RECT 242.4375 67.7700 242.7075 67.9950 ;
		LAYER VIA3 ;
        RECT 242.4375 67.7700 242.7075 67.9950 ;
		LAYER M2 ;
        RECT 242.4375 67.7700 242.7075 67.9950 ;
		LAYER M1 ;
        RECT 242.4375 77.3475 242.7075 77.4375 ;
		LAYER M3 ;
        RECT 242.4375 75.7800 242.7075 76.3275 ;
		LAYER VIA3 ;
        RECT 242.4375 75.7800 242.7075 76.3275 ;
		LAYER VIA3 ;
        RECT 242.4375 65.6250 242.7075 66.1200 ;
		LAYER M3 ;
        RECT 242.4375 64.9350 242.7075 65.1600 ;
		LAYER VIA3 ;
        RECT 242.4375 64.9350 242.7075 65.1600 ;
		LAYER M3 ;
        RECT 242.4375 62.7900 242.7075 63.2850 ;
		LAYER M3 ;
        RECT 242.4375 65.6250 242.7075 66.1200 ;
		LAYER M1 ;
        RECT 242.4375 62.0700 242.7075 62.3550 ;
		LAYER VIA3 ;
        RECT 242.4375 62.7900 242.7075 63.2850 ;
		LAYER VIA3 ;
        RECT 242.4375 62.1000 242.7075 62.3250 ;
		LAYER M3 ;
        RECT 242.4375 77.8725 242.7075 80.4150 ;
		LAYER VIA3 ;
        RECT 242.4375 77.8725 242.7075 80.4150 ;
		LAYER M2 ;
        RECT 242.4375 80.8800 242.7075 81.5850 ;
		LAYER M3 ;
        RECT 242.4375 80.8800 242.7075 81.5850 ;
		LAYER M2 ;
        RECT 242.4375 77.8725 242.7075 80.4150 ;
		LAYER VIA3 ;
        RECT 242.4375 80.8800 242.7075 81.5850 ;
		LAYER M3 ;
        RECT 242.4375 82.0500 242.7075 82.7175 ;
		LAYER M1 ;
        RECT 242.4375 82.0200 242.7075 82.7475 ;
		LAYER M2 ;
        RECT 242.4375 83.1825 242.7075 83.2125 ;
		LAYER M1 ;
        RECT 242.4375 83.1525 242.7075 83.2425 ;
		LAYER M2 ;
        RECT 242.4375 83.6775 242.7075 83.7075 ;
		LAYER M3 ;
        RECT 242.4375 83.6775 242.7075 83.7075 ;
		LAYER M3 ;
        RECT 242.4375 84.1725 242.7075 84.7125 ;
		LAYER VIA3 ;
        RECT 242.4375 84.1725 242.7075 84.7125 ;
		LAYER M1 ;
        RECT 242.4375 85.6425 242.7075 86.2350 ;
		LAYER M2 ;
        RECT 242.4375 85.1775 242.7075 85.2075 ;
		LAYER VIA3 ;
        RECT 242.4375 85.1775 242.7075 85.2075 ;
		LAYER M1 ;
        RECT 242.4375 84.1425 242.7075 84.7425 ;
		LAYER M1 ;
        RECT 242.4375 85.1475 242.7075 85.2375 ;
		LAYER M1 ;
        RECT 242.4375 86.6400 242.7075 87.2025 ;
		LAYER VIA3 ;
        RECT 242.4375 82.0500 242.7075 82.7175 ;
		LAYER M1 ;
        RECT 242.4375 91.5825 242.7075 91.7025 ;
		LAYER M1 ;
        RECT 242.4375 75.0600 242.7075 75.3450 ;
		LAYER M1 ;
        RECT 242.4375 111.0000 242.7075 111.5625 ;
		LAYER M3 ;
        RECT 242.4375 111.9975 242.7075 112.0275 ;
		LAYER VIA3 ;
        RECT 242.4375 111.9975 242.7075 112.0275 ;
		LAYER M2 ;
        RECT 242.4375 111.9975 242.7075 112.0275 ;
		LAYER M2 ;
        RECT 242.4375 75.7800 242.7075 76.3275 ;
		LAYER M1 ;
        RECT 242.4375 75.7500 242.7075 76.3575 ;
		LAYER M2 ;
        RECT 242.4375 76.7925 242.7075 76.9125 ;
		LAYER M1 ;
        RECT 242.4375 76.7625 242.7075 76.9425 ;
		LAYER M3 ;
        RECT 242.4375 76.7925 242.7075 76.9125 ;
		LAYER VIA3 ;
        RECT 242.4375 76.7925 242.7075 76.9125 ;
		LAYER M2 ;
        RECT 242.4375 68.4600 242.7075 68.9550 ;
		LAYER M2 ;
        RECT 242.4375 84.1725 242.7075 84.7125 ;
		LAYER M1 ;
        RECT 242.4375 80.8500 242.7075 81.6150 ;
		LAYER M1 ;
        RECT 242.4375 67.2450 242.7075 67.3350 ;
		LAYER M2 ;
        RECT 242.4375 59.9250 242.7075 60.4500 ;
		LAYER M3 ;
        RECT 242.4375 59.9250 242.7075 60.4500 ;
		LAYER M3 ;
        RECT 242.4375 61.6050 242.7075 61.6350 ;
		LAYER M2 ;
        RECT 242.4375 60.9150 242.7075 61.1400 ;
		LAYER M3 ;
        RECT 242.4375 60.9150 242.7075 61.1400 ;
		LAYER M1 ;
        RECT 242.4375 60.8850 242.7075 61.1700 ;
		LAYER M3 ;
        RECT 242.4375 88.1325 242.7075 88.1925 ;
		LAYER M1 ;
        RECT 242.4375 88.1025 242.7075 88.2225 ;
		LAYER M2 ;
        RECT 242.4375 87.6375 242.7075 87.6675 ;
		LAYER M3 ;
        RECT 242.4375 87.6375 242.7075 87.6675 ;
		LAYER M3 ;
        RECT 242.4375 88.6575 242.7075 88.6875 ;
		LAYER M3 ;
        RECT 242.4375 91.1175 242.7075 91.1475 ;
		LAYER M2 ;
        RECT 242.4375 91.1175 242.7075 91.1475 ;
		LAYER VIA3 ;
        RECT 242.4375 88.6575 242.7075 88.6875 ;
		LAYER M1 ;
        RECT 242.4375 89.1225 242.7075 89.7150 ;
		LAYER M2 ;
        RECT 242.4375 88.6575 242.7075 88.6875 ;
		LAYER VIA3 ;
        RECT 242.4375 91.1175 242.7075 91.1475 ;
		LAYER VIA3 ;
        RECT 242.4375 86.6700 242.7075 87.1725 ;
		LAYER M2 ;
        RECT 242.4375 86.6700 242.7075 87.1725 ;
		LAYER M1 ;
        RECT 242.4375 87.6075 242.7075 87.6975 ;
		LAYER M3 ;
        RECT 242.4375 86.6700 242.7075 87.1725 ;
		LAYER M1 ;
        RECT 242.4375 88.6275 242.7075 88.7175 ;
		LAYER M2 ;
        RECT 242.4375 89.1525 242.7075 89.6850 ;
		LAYER M3 ;
        RECT 242.4375 89.1525 242.7075 89.6850 ;
		LAYER VIA3 ;
        RECT 242.4375 89.1525 242.7075 89.6850 ;
		LAYER VIA3 ;
        RECT 242.4375 90.1500 242.7075 90.6525 ;
		LAYER M2 ;
        RECT 242.4375 90.1500 242.7075 90.6525 ;
		LAYER M3 ;
        RECT 242.4375 90.1500 242.7075 90.6525 ;
		LAYER M1 ;
        RECT 242.4375 90.1200 242.7075 90.6825 ;
		LAYER VIA3 ;
        RECT 242.4375 88.1325 242.7075 88.1925 ;
		LAYER M2 ;
        RECT 242.4375 88.1325 242.7075 88.1925 ;
		LAYER VIA3 ;
        RECT 242.4375 87.6375 242.7075 87.6675 ;
		LAYER M2 ;
        RECT 242.4375 99.0975 242.7075 99.1275 ;
		LAYER M2 ;
        RECT 242.4375 95.6175 242.7075 95.6475 ;
		LAYER M1 ;
        RECT 242.4375 95.5875 242.7075 95.6775 ;
		LAYER VIA3 ;
        RECT 242.4375 99.0975 242.7075 99.1275 ;
		LAYER M3 ;
        RECT 242.4375 95.0925 242.7075 95.1525 ;
		LAYER VIA3 ;
        RECT 242.4375 95.0925 242.7075 95.1525 ;
		LAYER M1 ;
        RECT 242.4375 95.0625 242.7075 95.1825 ;
		LAYER M3 ;
        RECT 242.4375 95.6175 242.7075 95.6475 ;
		LAYER M2 ;
        RECT 242.4375 95.0925 242.7075 95.1525 ;
		LAYER VIA3 ;
        RECT 242.4375 95.6175 242.7075 95.6475 ;
		LAYER VIA3 ;
        RECT 242.4375 94.5975 242.7075 94.6275 ;
		LAYER M1 ;
        RECT 242.4375 94.5675 242.7075 94.6575 ;
		LAYER M2 ;
        RECT 242.4375 93.6300 242.7075 94.1325 ;
		LAYER VIA3 ;
        RECT 242.4375 93.6300 242.7075 94.1325 ;
		LAYER M3 ;
        RECT 242.4375 94.5975 242.7075 94.6275 ;
		LAYER M2 ;
        RECT 242.4375 94.5975 242.7075 94.6275 ;
		LAYER M2 ;
        RECT 242.4375 98.0775 242.7075 98.1075 ;
		LAYER M3 ;
        RECT 242.4375 96.1125 242.7075 96.6450 ;
		LAYER VIA3 ;
        RECT 242.4375 96.1125 242.7075 96.6450 ;
		LAYER M2 ;
        RECT 242.4375 96.1125 242.7075 96.6450 ;
		LAYER M2 ;
        RECT 242.4375 91.6125 242.7075 91.6725 ;
		LAYER M3 ;
        RECT 242.4375 91.6125 242.7075 91.6725 ;
		LAYER VIA3 ;
        RECT 242.4375 91.6125 242.7075 91.6725 ;
		LAYER M1 ;
        RECT 242.4375 99.0675 242.7075 99.1575 ;
		LAYER M1 ;
        RECT 242.4375 101.5275 242.7075 101.6175 ;
		LAYER M3 ;
        RECT 242.4375 101.5575 242.7075 101.5875 ;
		LAYER VIA3 ;
        RECT 242.4375 101.5575 242.7075 101.5875 ;
		LAYER M2 ;
        RECT 242.4375 101.5575 242.7075 101.5875 ;
		LAYER M1 ;
        RECT 242.4375 100.5600 242.7075 101.1225 ;
		LAYER M2 ;
        RECT 242.4375 92.1375 242.7075 92.1675 ;
		LAYER M3 ;
        RECT 242.4375 92.1375 242.7075 92.1675 ;
		LAYER VIA3 ;
        RECT 242.4375 92.1375 242.7075 92.1675 ;
		LAYER M1 ;
        RECT 242.4375 92.1075 242.7075 92.1975 ;
		LAYER M2 ;
        RECT 242.4375 92.6325 242.7075 93.1650 ;
		LAYER M3 ;
        RECT 242.4375 92.6325 242.7075 93.1650 ;
		LAYER M1 ;
        RECT 242.4375 92.6025 242.7075 93.1950 ;
		LAYER M1 ;
        RECT 242.4375 93.6000 242.7075 94.1625 ;
		LAYER M3 ;
        RECT 242.4375 99.0975 242.7075 99.1275 ;
		LAYER M2 ;
        RECT 242.4375 102.0525 242.7075 102.1125 ;
		LAYER M1 ;
        RECT 242.4375 102.0225 242.7075 102.1425 ;
		LAYER M3 ;
        RECT 242.4375 102.0525 242.7075 102.1125 ;
		LAYER M3 ;
        RECT 242.4375 103.0725 242.7075 103.6050 ;
		LAYER VIA3 ;
        RECT 242.4375 103.0725 242.7075 103.6050 ;
		LAYER M3 ;
        RECT 242.4375 102.5775 242.7075 102.6075 ;
		LAYER VIA3 ;
        RECT 242.4375 102.5775 242.7075 102.6075 ;
		LAYER VIA3 ;
        RECT 242.4375 77.3775 242.7075 77.4075 ;
		LAYER M2 ;
        RECT 242.4375 77.3775 242.7075 77.4075 ;
		LAYER M3 ;
        RECT 242.4375 77.3775 242.7075 77.4075 ;
		LAYER VIA3 ;
        RECT 242.4375 85.6725 242.7075 86.2050 ;
		LAYER M1 ;
        RECT 242.4375 83.6475 242.7075 83.7375 ;
		LAYER M3 ;
        RECT 242.4375 83.1825 242.7075 83.2125 ;
		LAYER M2 ;
        RECT 242.4375 82.0500 242.7075 82.7175 ;
		LAYER VIA3 ;
        RECT 242.4375 83.1825 242.7075 83.2125 ;
		LAYER M2 ;
        RECT 242.4375 85.6725 242.7075 86.2050 ;
		LAYER M3 ;
        RECT 242.4375 85.6725 242.7075 86.2050 ;
		LAYER M1 ;
        RECT 242.4375 91.0875 242.7075 91.1775 ;
		LAYER M3 ;
        RECT 242.4375 107.5500 242.7075 108.0525 ;
		LAYER VIA3 ;
        RECT 242.4375 105.5325 242.7075 105.5925 ;
		LAYER M2 ;
        RECT 242.4375 106.5525 242.7075 107.0850 ;
		LAYER M2 ;
        RECT 242.4375 108.5175 242.7075 108.5475 ;
		LAYER M2 ;
        RECT 242.4375 107.5500 242.7075 108.0525 ;
		LAYER M1 ;
        RECT 242.4375 108.4875 242.7075 108.5775 ;
		LAYER M3 ;
        RECT 242.4375 108.5175 242.7075 108.5475 ;
		LAYER VIA3 ;
        RECT 242.4375 108.5175 242.7075 108.5475 ;
		LAYER VIA3 ;
        RECT 242.4375 107.5500 242.7075 108.0525 ;
		LAYER M1 ;
        RECT 242.4375 104.0400 242.7075 104.6025 ;
		LAYER M3 ;
        RECT 242.4375 105.5325 242.7075 105.5925 ;
		LAYER M1 ;
        RECT 242.4375 105.0075 242.7075 105.0975 ;
		LAYER VIA3 ;
        RECT 242.4375 104.0700 242.7075 104.5725 ;
		LAYER M3 ;
        RECT 242.4375 109.5375 242.7075 109.5675 ;
		LAYER VIA3 ;
        RECT 242.4375 110.0325 242.7075 110.5650 ;
		LAYER M1 ;
        RECT 242.4375 110.0025 242.7075 110.5950 ;
		LAYER M1 ;
        RECT 242.4375 107.5200 242.7075 108.0825 ;
		LAYER VIA3 ;
        RECT 242.4375 109.5375 242.7075 109.5675 ;
		LAYER M1 ;
        RECT 242.4375 109.5075 242.7075 109.5975 ;
		LAYER VIA3 ;
        RECT 242.4375 106.0575 242.7075 106.0875 ;
		LAYER M2 ;
        RECT 242.4375 106.0575 242.7075 106.0875 ;
		LAYER M1 ;
        RECT 242.4375 106.0275 242.7075 106.1175 ;
		LAYER M2 ;
        RECT 242.4375 105.5325 242.7075 105.5925 ;
		LAYER M3 ;
        RECT 242.4375 109.0125 242.7075 109.0725 ;
		LAYER M2 ;
        RECT 242.4375 109.0125 242.7075 109.0725 ;
		LAYER VIA3 ;
        RECT 242.4375 109.0125 242.7075 109.0725 ;
		LAYER M1 ;
        RECT 242.4375 108.9825 242.7075 109.1025 ;
		LAYER M3 ;
        RECT 242.4375 98.0775 242.7075 98.1075 ;
		LAYER VIA3 ;
        RECT 242.4375 98.0775 242.7075 98.1075 ;
		LAYER M1 ;
        RECT 242.4375 96.0825 242.7075 96.6750 ;
		LAYER M3 ;
        RECT 242.4375 97.1100 242.7075 97.6125 ;
		LAYER M2 ;
        RECT 242.4375 97.1100 242.7075 97.6125 ;
		LAYER VIA3 ;
        RECT 242.4375 99.5925 242.7075 100.1250 ;
		LAYER M2 ;
        RECT 242.4375 99.5925 242.7075 100.1250 ;
		LAYER M3 ;
        RECT 242.4375 99.5925 242.7075 100.1250 ;
		LAYER M1 ;
        RECT 242.4375 99.5625 242.7075 100.1550 ;
		LAYER M2 ;
        RECT 242.4375 100.5900 242.7075 101.0925 ;
		LAYER M3 ;
        RECT 242.4375 100.5900 242.7075 101.0925 ;
		LAYER VIA3 ;
        RECT 242.4375 100.5900 242.7075 101.0925 ;
		LAYER M1 ;
        RECT 242.4375 140.3025 242.7075 141.6150 ;
		LAYER M2 ;
        RECT 242.4375 140.3325 242.7075 141.6150 ;
		LAYER VIA3 ;
        RECT 242.4375 140.3325 242.7075 141.6150 ;
		LAYER M1 ;
        RECT 242.4375 133.8675 242.7075 133.9575 ;
		LAYER M3 ;
        RECT 242.4375 139.8375 242.7075 139.8675 ;
		LAYER M3 ;
        RECT 242.4375 120.4725 242.7075 121.0050 ;
		LAYER VIA3 ;
        RECT 242.4375 120.4725 242.7075 121.0050 ;
		LAYER M2 ;
        RECT 242.4375 121.4700 242.7075 121.9725 ;
		LAYER M3 ;
        RECT 242.4375 106.0575 242.7075 106.0875 ;
		LAYER M3 ;
        RECT 242.4375 106.5525 242.7075 107.0850 ;
		LAYER VIA3 ;
        RECT 242.4375 106.5525 242.7075 107.0850 ;
		LAYER M1 ;
        RECT 242.4375 98.0475 242.7075 98.1375 ;
		LAYER VIA3 ;
        RECT 242.4375 98.5725 242.7075 98.6325 ;
		LAYER M3 ;
        RECT 242.4375 98.5725 242.7075 98.6325 ;
		LAYER M2 ;
        RECT 242.4375 98.5725 242.7075 98.6325 ;
		LAYER M3 ;
        RECT 242.4375 140.3325 242.7075 141.6150 ;
		LAYER M3 ;
        RECT 242.4375 133.3725 242.7075 133.4325 ;
		LAYER VIA3 ;
        RECT 242.4375 133.3725 242.7075 133.4325 ;
		LAYER M1 ;
        RECT 242.4375 137.3475 242.7075 137.4375 ;
		LAYER VIA3 ;
        RECT 242.4375 136.8525 242.7075 136.9125 ;
		LAYER VIA3 ;
        RECT 242.4375 136.3575 242.7075 136.3875 ;
		LAYER M2 ;
        RECT 242.4375 134.3925 242.7075 134.9250 ;
		LAYER VIA3 ;
        RECT 242.4375 131.9100 242.7075 132.4125 ;
		LAYER M2 ;
        RECT 242.4375 128.4300 242.7075 128.9325 ;
		LAYER M1 ;
        RECT 242.4375 127.4025 242.7075 127.9950 ;
		LAYER M2 ;
        RECT 242.4375 130.4175 242.7075 130.4475 ;
		LAYER M1 ;
        RECT 242.4375 134.3625 242.7075 134.9550 ;
		LAYER M3 ;
        RECT 242.4375 126.9375 242.7075 126.9675 ;
		LAYER M1 ;
        RECT 242.4375 126.9075 242.7075 126.9975 ;
		LAYER M2 ;
        RECT 242.4375 133.3725 242.7075 133.4325 ;
		LAYER M4 ;
        RECT 0.0000 95.6325 242.1300 98.0925 ;
		LAYER M4 ;
        RECT 0.0000 99.1125 242.1300 101.5725 ;
		LAYER M4 ;
        RECT 0.0000 102.5925 242.1300 105.0525 ;
		LAYER M4 ;
        RECT 0.0000 5.2425 242.1300 7.7025 ;
		LAYER M4 ;
        RECT 0.0000 1.7625 242.1300 4.2225 ;
		LAYER VIA2 ;
        RECT 0.0000 0.0000 242.7075 141.6150 ;
		LAYER M4 ;
        RECT 0.0000 58.9350 106.9050 59.6325 ;
		LAYER M4 ;
        RECT 0.0000 0.0000 242.1300 1.1775 ;
		LAYER M4 ;
        RECT 0.0000 40.0425 242.1300 42.5025 ;
		LAYER M4 ;
        RECT 0.0000 50.4825 242.1300 52.9425 ;
		LAYER M4 ;
        RECT 0.0000 92.1525 242.1300 94.6125 ;
		LAYER M3 ;
        RECT 0.0000 0.0000 242.4375 141.6150 ;
		LAYER M2 ;
        RECT 0.0000 0.0000 242.4375 141.6150 ;
		LAYER VIA3 ;
        RECT 0.0000 0.0000 242.4375 141.6150 ;
		LAYER M4 ;
        RECT 0.0000 22.6425 242.1300 25.1025 ;
		LAYER M4 ;
        RECT 0.0000 19.1625 242.1300 21.6225 ;
		LAYER M4 ;
        RECT 0.0000 12.2025 242.1300 14.6625 ;
		LAYER M4 ;
        RECT 0.0000 8.7225 242.1300 11.1825 ;
		LAYER M2 ;
        RECT 242.4375 69.4200 242.7075 69.6450 ;
		LAYER M4 ;
        RECT 0.0000 68.8050 242.2050 72.6075 ;
		LAYER M4 ;
        RECT 0.0000 65.1675 242.2050 68.1750 ;
		LAYER M4 ;
        RECT 0.0000 78.3225 242.2050 80.9250 ;
		LAYER M4 ;
        RECT 0.0000 73.2375 242.2050 75.6375 ;
		LAYER M4 ;
        RECT 0.0000 76.2675 242.2050 77.6925 ;
		LAYER M4 ;
        RECT 106.9050 56.9325 132.5100 59.6325 ;
		LAYER M4 ;
        RECT 132.5100 58.9350 238.1400 59.6325 ;
		LAYER M4 ;
        RECT 0.0000 57.0075 242.1300 59.4825 ;
		LAYER M4 ;
        RECT 0.0000 60.2625 242.2050 62.0025 ;
		LAYER M4 ;
        RECT 0.0000 53.9625 242.1300 56.4225 ;
		LAYER M4 ;
        RECT 0.0000 62.6325 242.2050 64.5375 ;
		LAYER M4 ;
        RECT 0.0000 85.1925 242.1300 87.6525 ;
		LAYER M4 ;
        RECT 0.0000 88.6725 242.1300 91.1325 ;
		LAYER M4 ;
        RECT 0.0000 81.5550 242.2050 84.6825 ;
		LAYER M4 ;
        RECT 0.0000 130.4325 242.1300 132.8925 ;
		LAYER M4 ;
        RECT 0.0000 133.9125 242.1300 136.3725 ;
		LAYER M4 ;
        RECT 0.0000 137.3925 242.1300 139.8525 ;
		LAYER M4 ;
        RECT 0.0000 140.4375 242.1300 141.6150 ;
		LAYER M4 ;
        RECT 0.0000 113.0325 242.1300 115.4925 ;
		LAYER M4 ;
        RECT 0.0000 109.5525 242.1300 112.0125 ;
		LAYER M4 ;
        RECT 0.0000 106.0725 242.1300 108.5325 ;
		LAYER M4 ;
        RECT 0.0000 116.5125 242.1300 118.9725 ;
		LAYER M4 ;
        RECT 0.0000 119.9925 242.1300 122.4525 ;
		LAYER M4 ;
        RECT 0.0000 123.4725 242.1300 125.9325 ;
		LAYER M4 ;
        RECT 0.0000 126.9525 242.1300 129.4125 ;
		LAYER M4 ;
        RECT 0.0000 43.5225 242.1300 45.9825 ;
		LAYER M4 ;
        RECT 0.0000 47.0025 242.1300 49.4625 ;
		LAYER M4 ;
        RECT 0.0000 36.5625 242.1300 39.0225 ;
		LAYER M4 ;
        RECT 0.0000 33.0825 242.1300 35.5425 ;
		LAYER M4 ;
        RECT 0.0000 29.6025 242.1300 32.0625 ;
		LAYER M4 ;
        RECT 0.0000 15.6825 242.1300 18.1425 ;
		LAYER M4 ;
        RECT 0.0000 26.1225 242.1300 28.5825 ;
		LAYER M4 ;
        RECT 242.1300 0.0000 242.2050 59.4825 ;
		LAYER VIA1 ;
        RECT 0.0000 0.0000 242.7075 141.6150 ;
		LAYER M1 ;
        RECT 0.0000 0.0000 242.4375 141.6150 ;
		LAYER M1 ;
        RECT 242.4375 139.8075 242.7075 139.8975 ;
		LAYER M2 ;
        RECT 242.4375 66.5850 242.7075 66.8100 ;
		LAYER M1 ;
        RECT 242.4375 65.5950 242.7075 66.1500 ;
		LAYER M2 ;
        RECT 242.4375 138.8700 242.7075 139.3725 ;
		LAYER M1 ;
        RECT 242.4375 138.8400 242.7075 139.4025 ;
		LAYER M2 ;
        RECT 242.4375 137.3775 242.7075 137.4075 ;
		LAYER M3 ;
        RECT 242.4375 68.4600 242.7075 68.9550 ;
		LAYER M3 ;
        RECT 242.4375 69.4200 242.7075 69.6450 ;
		LAYER M1 ;
        RECT 242.4375 9.1725 242.7075 9.7650 ;
		LAYER M2 ;
        RECT 242.4375 9.2025 242.7075 9.7350 ;
		LAYER M3 ;
        RECT 242.4375 10.2000 242.7075 10.7025 ;
		LAYER M1 ;
        RECT 242.4375 10.1700 242.7075 10.7325 ;
		LAYER M4 ;
        RECT 238.1400 56.9325 239.4000 59.6325 ;
		LAYER M2 ;
        RECT 242.4375 11.1675 242.7075 11.1975 ;
		LAYER M4 ;
        RECT 239.4000 58.9350 242.2050 59.6325 ;
		LAYER M2 ;
        RECT 242.4375 15.6675 242.7075 15.6975 ;
		LAYER M2 ;
        RECT 242.4375 14.6475 242.7075 14.6775 ;
		LAYER M3 ;
        RECT 242.4375 14.6475 242.7075 14.6775 ;
		LAYER M1 ;
        RECT 242.4375 14.6175 242.7075 14.7075 ;
		LAYER VIA3 ;
        RECT 242.4375 15.6675 242.7075 15.6975 ;
		LAYER M2 ;
        RECT 242.4375 54.4425 242.7075 54.9750 ;
		LAYER M1 ;
        RECT 242.4375 54.4125 242.7075 55.0050 ;
		LAYER VIA3 ;
        RECT 242.4375 53.9475 242.7075 53.9775 ;
		LAYER M2 ;
        RECT 242.4375 53.9475 242.7075 53.9775 ;
		LAYER VIA3 ;
        RECT 242.4375 54.4425 242.7075 54.9750 ;
		LAYER M1 ;
        RECT 242.4375 48.4500 242.7075 49.0125 ;
		LAYER VIA3 ;
        RECT 242.4375 47.4825 242.7075 48.0150 ;
		LAYER M1 ;
        RECT 242.4375 47.4525 242.7075 48.0450 ;
		LAYER VIA3 ;
        RECT 242.4375 46.9875 242.7075 47.0175 ;
		LAYER M1 ;
        RECT 242.4375 77.8425 242.7075 80.4450 ;
		LAYER M2 ;
        RECT 242.4375 70.1100 242.7075 70.1400 ;
		LAYER M3 ;
        RECT 242.4375 70.1100 242.7075 70.1400 ;
		LAYER M4 ;
        RECT 242.1300 81.7050 242.2050 141.6150 ;
		LAYER M3 ;
        RECT 242.4375 123.4575 242.7075 123.4875 ;
		LAYER VIA3 ;
        RECT 242.4375 123.4575 242.7075 123.4875 ;
		LAYER M1 ;
        RECT 242.4375 123.4275 242.7075 123.5175 ;
		LAYER M3 ;
        RECT 242.4375 85.1775 242.7075 85.2075 ;
		LAYER VIA3 ;
        RECT 242.4375 83.6775 242.7075 83.7075 ;
		LAYER M1 ;
        RECT 242.4375 97.0800 242.7075 97.6425 ;
		LAYER M1 ;
        RECT 242.4375 122.9025 242.7075 123.0225 ;
		LAYER M2 ;
        RECT 242.4375 123.4575 242.7075 123.4875 ;
		LAYER M1 ;
        RECT 242.4375 106.5225 242.7075 107.1150 ;
		LAYER VIA3 ;
        RECT 242.4375 97.1100 242.7075 97.6125 ;
		LAYER M1 ;
        RECT 242.4375 98.5425 242.7075 98.6625 ;
		LAYER M1 ;
        RECT 242.4375 74.1000 242.7075 74.6550 ;
		LAYER M1 ;
        RECT 242.4375 72.9150 242.7075 73.0050 ;
		LAYER M2 ;
        RECT 242.4375 72.2550 242.7075 72.4800 ;
		LAYER VIA3 ;
        RECT 242.4375 70.1100 242.7075 70.1400 ;
		LAYER M3 ;
        RECT 242.4375 72.9450 242.7075 72.9750 ;
		LAYER M3 ;
        RECT 242.4375 11.1675 242.7075 11.1975 ;
		LAYER M2 ;
        RECT 242.4375 8.1825 242.7075 8.2425 ;
		LAYER M3 ;
        RECT 242.4375 8.1825 242.7075 8.2425 ;
		LAYER M1 ;
        RECT 242.4375 11.1375 242.7075 11.2275 ;
		LAYER M2 ;
        RECT 242.4375 10.2000 242.7075 10.7025 ;
		LAYER M1 ;
        RECT 242.4375 11.6325 242.7075 11.7525 ;
		LAYER VIA3 ;
        RECT 242.4375 11.1675 242.7075 11.1975 ;
		LAYER VIA3 ;
        RECT 242.4375 10.2000 242.7075 10.7025 ;
		LAYER VIA3 ;
        RECT 242.4375 42.9825 242.7075 43.0425 ;
		LAYER M3 ;
        RECT 242.4375 42.9825 242.7075 43.0425 ;
		LAYER M1 ;
        RECT 242.4375 42.9525 242.7075 43.0725 ;
		LAYER VIA3 ;
        RECT 242.4375 42.4875 242.7075 42.5175 ;
		LAYER M3 ;
        RECT 242.4375 42.4875 242.7075 42.5175 ;
		LAYER VIA3 ;
        RECT 242.4375 41.5200 242.7075 42.0225 ;
		LAYER M1 ;
        RECT 242.4375 44.9700 242.7075 45.5325 ;
		LAYER M2 ;
        RECT 242.4375 42.4875 242.7075 42.5175 ;
		LAYER M3 ;
        RECT 242.4375 9.2025 242.7075 9.7350 ;
		LAYER VIA3 ;
        RECT 242.4375 8.7075 242.7075 8.7375 ;
		LAYER M3 ;
        RECT 242.4375 8.7075 242.7075 8.7375 ;
		LAYER M1 ;
        RECT 242.4375 8.6775 242.7075 8.7675 ;
		LAYER VIA3 ;
        RECT 242.4375 9.2025 242.7075 9.7350 ;
		LAYER M2 ;
        RECT 242.4375 8.7075 242.7075 8.7375 ;
		LAYER VIA3 ;
        RECT 242.4375 7.6875 242.7075 7.7175 ;
		LAYER M2 ;
        RECT 242.4375 7.6875 242.7075 7.7175 ;
		LAYER M3 ;
        RECT 242.4375 7.6875 242.7075 7.7175 ;
		LAYER VIA3 ;
        RECT 242.4375 8.1825 242.7075 8.2425 ;
		LAYER M1 ;
        RECT 242.4375 8.1525 242.7075 8.2725 ;
		LAYER M1 ;
        RECT 242.4375 46.9575 242.7075 47.0475 ;
		LAYER M1 ;
        RECT 242.4375 45.9375 242.7075 46.0275 ;
		LAYER VIA3 ;
        RECT 242.4375 45.9675 242.7075 45.9975 ;
		LAYER VIA3 ;
        RECT 242.4375 46.4625 242.7075 46.5225 ;
		LAYER M2 ;
        RECT 242.4375 46.4625 242.7075 46.5225 ;
		LAYER M1 ;
        RECT 242.4375 46.4325 242.7075 46.5525 ;
		LAYER M3 ;
        RECT 242.4375 45.9675 242.7075 45.9975 ;
		LAYER VIA3 ;
        RECT 242.4375 45.0000 242.7075 45.5025 ;
		LAYER M2 ;
        RECT 242.4375 45.0000 242.7075 45.5025 ;
		LAYER M3 ;
        RECT 242.4375 44.0025 242.7075 44.5350 ;
		LAYER M3 ;
        RECT 242.4375 45.0000 242.7075 45.5025 ;
		LAYER VIA3 ;
        RECT 242.4375 43.5075 242.7075 43.5375 ;
		LAYER M2 ;
        RECT 242.4375 43.5075 242.7075 43.5375 ;
		LAYER M1 ;
        RECT 242.4375 43.4775 242.7075 43.5675 ;
		LAYER M2 ;
        RECT 242.4375 44.0025 242.7075 44.5350 ;
		LAYER M1 ;
        RECT 242.4375 43.9725 242.7075 44.5650 ;
		LAYER M2 ;
        RECT 242.4375 1.7475 242.7075 1.7775 ;
		LAYER M3 ;
        RECT 242.4375 3.2400 242.7075 3.7425 ;
		LAYER VIA3 ;
        RECT 242.4375 3.2400 242.7075 3.7425 ;
		LAYER M2 ;
        RECT 242.4375 5.2275 242.7075 5.2575 ;
		LAYER VIA3 ;
        RECT 242.4375 5.2275 242.7075 5.2575 ;
		LAYER VIA3 ;
        RECT 242.4375 4.7025 242.7075 4.7625 ;
		LAYER M2 ;
        RECT 242.4375 4.7025 242.7075 4.7625 ;
		LAYER M3 ;
        RECT 242.4375 4.7025 242.7075 4.7625 ;
		LAYER M3 ;
        RECT 242.4375 5.2275 242.7075 5.2575 ;
		LAYER M2 ;
        RECT 242.4375 5.7225 242.7075 6.2550 ;
		LAYER M3 ;
        RECT 242.4375 5.7225 242.7075 6.2550 ;
		LAYER M1 ;
        RECT 242.4375 5.1975 242.7075 5.2875 ;
		LAYER M1 ;
        RECT 242.4375 4.6725 242.7075 4.7925 ;
		LAYER VIA3 ;
        RECT 242.4375 5.7225 242.7075 6.2550 ;
		LAYER VIA3 ;
        RECT 242.4375 4.2075 242.7075 4.2375 ;
		LAYER M2 ;
        RECT 242.4375 6.7200 242.7075 7.2225 ;
		LAYER M3 ;
        RECT 242.4375 6.7200 242.7075 7.2225 ;
		LAYER M1 ;
        RECT 242.4375 5.6925 242.7075 6.2850 ;
		LAYER M1 ;
        RECT 242.4375 4.1775 242.7075 4.2675 ;
		LAYER VIA3 ;
        RECT 242.4375 6.7200 242.7075 7.2225 ;
		LAYER M2 ;
        RECT 242.4375 2.2425 242.7075 2.7750 ;
		LAYER M3 ;
        RECT 242.4375 2.2425 242.7075 2.7750 ;
		LAYER VIA3 ;
        RECT 242.4375 2.2425 242.7075 2.7750 ;
		LAYER M2 ;
        RECT 242.4375 3.2400 242.7075 3.7425 ;
		LAYER M1 ;
        RECT 242.4375 3.2100 242.7075 3.7725 ;
		LAYER M1 ;
        RECT 242.4375 53.9175 242.7075 54.0075 ;
		LAYER M2 ;
        RECT 242.4375 53.4225 242.7075 53.4825 ;
		LAYER M3 ;
        RECT 242.4375 53.4225 242.7075 53.4825 ;
		LAYER M2 ;
        RECT 242.4375 49.4475 242.7075 49.4775 ;
		LAYER VIA3 ;
        RECT 242.4375 49.4475 242.7075 49.4775 ;
		LAYER M3 ;
        RECT 242.4375 49.9425 242.7075 50.0025 ;
		LAYER M2 ;
        RECT 242.4375 48.4800 242.7075 48.9825 ;
		LAYER M1 ;
        RECT 242.4375 7.6575 242.7075 7.7475 ;
		LAYER M1 ;
        RECT 242.4375 6.6900 242.7075 7.2525 ;
		LAYER M3 ;
        RECT 242.4375 48.4800 242.7075 48.9825 ;
		LAYER M2 ;
        RECT 242.4375 4.2075 242.7075 4.2375 ;
		LAYER M3 ;
        RECT 242.4375 4.2075 242.7075 4.2375 ;
		LAYER M1 ;
        RECT 242.4375 64.4100 242.7075 64.5000 ;
		LAYER M2 ;
        RECT 242.4375 64.4400 242.7075 64.4700 ;
		LAYER M3 ;
        RECT 242.4375 64.4400 242.7075 64.4700 ;
		LAYER M2 ;
        RECT 242.4375 64.9350 242.7075 65.1600 ;
		LAYER VIA3 ;
        RECT 242.4375 64.4400 242.7075 64.4700 ;
		LAYER M2 ;
        RECT 242.4375 65.6250 242.7075 66.1200 ;
		LAYER VIA3 ;
        RECT 242.4375 66.5850 242.7075 66.8100 ;
		LAYER M1 ;
        RECT 242.4375 64.9050 242.7075 65.1900 ;
		LAYER M2 ;
        RECT 242.4375 63.7500 242.7075 63.9750 ;
		LAYER VIA3 ;
        RECT 242.4375 63.7500 242.7075 63.9750 ;
		LAYER M1 ;
        RECT 242.4375 63.7200 242.7075 64.0050 ;
		LAYER M2 ;
        RECT 242.4375 62.7900 242.7075 63.2850 ;
		LAYER M1 ;
        RECT 242.4375 62.7600 242.7075 63.3150 ;
		LAYER M2 ;
        RECT 242.4375 61.6050 242.7075 61.6350 ;
		LAYER VIA3 ;
        RECT 242.4375 61.6050 242.7075 61.6350 ;
		LAYER M1 ;
        RECT 242.4375 61.5750 242.7075 61.6650 ;
		LAYER VIA3 ;
        RECT 242.4375 60.9150 242.7075 61.1400 ;
		LAYER M3 ;
        RECT 242.4375 133.8975 242.7075 133.9275 ;
		LAYER VIA3 ;
        RECT 242.4375 133.8975 242.7075 133.9275 ;
		LAYER M3 ;
        RECT 242.4375 131.9100 242.7075 132.4125 ;
		LAYER M1 ;
        RECT 242.4375 133.3425 242.7075 133.4625 ;
		LAYER M1 ;
        RECT 242.4375 105.5025 242.7075 105.6225 ;
		LAYER M2 ;
        RECT 242.4375 110.0325 242.7075 110.5650 ;
		LAYER M2 ;
        RECT 242.4375 111.0300 242.7075 111.5325 ;
		LAYER M3 ;
        RECT 242.4375 111.0300 242.7075 111.5325 ;
		LAYER M3 ;
        RECT 242.4375 110.0325 242.7075 110.5650 ;
		LAYER M2 ;
        RECT 242.4375 109.5375 242.7075 109.5675 ;
		LAYER M2 ;
        RECT 242.4375 104.0700 242.7075 104.5725 ;
		LAYER M3 ;
        RECT 242.4375 104.0700 242.7075 104.5725 ;
		LAYER VIA3 ;
        RECT 242.4375 111.0300 242.7075 111.5325 ;
		LAYER M3 ;
        RECT 242.4375 105.0375 242.7075 105.0675 ;
		LAYER M2 ;
        RECT 242.4375 105.0375 242.7075 105.0675 ;
		LAYER VIA3 ;
        RECT 242.4375 105.0375 242.7075 105.0675 ;
		LAYER M2 ;
        RECT 242.4375 133.8975 242.7075 133.9275 ;
		LAYER M1 ;
        RECT 242.4375 131.8800 242.7075 132.4425 ;
		LAYER M1 ;
        RECT 242.4375 130.3875 242.7075 130.4775 ;
		LAYER M3 ;
        RECT 242.4375 132.8775 242.7075 132.9075 ;
		LAYER M2 ;
        RECT 242.4375 132.8775 242.7075 132.9075 ;
		LAYER VIA3 ;
        RECT 242.4375 132.8775 242.7075 132.9075 ;
		LAYER M2 ;
        RECT 242.4375 131.9100 242.7075 132.4125 ;
		LAYER M2 ;
        RECT 242.4375 130.9125 242.7075 131.4450 ;
		LAYER VIA3 ;
        RECT 242.4375 130.9125 242.7075 131.4450 ;
		LAYER M3 ;
        RECT 242.4375 130.9125 242.7075 131.4450 ;
		LAYER M1 ;
        RECT 242.4375 130.8825 242.7075 131.4750 ;
		LAYER M2 ;
        RECT 242.4375 119.4525 242.7075 119.5125 ;
		LAYER M3 ;
        RECT 242.4375 119.4525 242.7075 119.5125 ;
		LAYER M1 ;
        RECT 242.4375 125.8875 242.7075 125.9775 ;
		LAYER M1 ;
        RECT 242.4375 102.5475 242.7075 102.6375 ;
		LAYER M3 ;
        RECT 242.4375 117.9900 242.7075 118.4925 ;
		LAYER M2 ;
        RECT 242.4375 118.9575 242.7075 118.9875 ;
		LAYER M1 ;
        RECT 242.4375 103.0425 242.7075 103.6350 ;
		LAYER M2 ;
        RECT 242.4375 103.0725 242.7075 103.6050 ;
		LAYER M2 ;
        RECT 242.4375 102.5775 242.7075 102.6075 ;
		LAYER VIA3 ;
        RECT 242.4375 102.0525 242.7075 102.1125 ;
		LAYER VIA3 ;
        RECT 242.4375 92.6325 242.7075 93.1650 ;
		LAYER M3 ;
        RECT 242.4375 93.6300 242.7075 94.1325 ;
		LAYER M1 ;
        RECT 242.4375 66.5550 242.7075 66.8400 ;
		LAYER M2 ;
        RECT 242.4375 67.2750 242.7075 67.3050 ;
		LAYER VIA3 ;
        RECT 242.4375 67.2750 242.7075 67.3050 ;
		LAYER M3 ;
        RECT 242.4375 67.2750 242.7075 67.3050 ;
		LAYER M3 ;
        RECT 242.4375 66.5850 242.7075 66.8100 ;
		LAYER M2 ;
        RECT 242.4375 62.1000 242.7075 62.3250 ;
		LAYER VIA3 ;
        RECT 242.4375 59.9250 242.7075 60.4500 ;
		LAYER M1 ;
        RECT 242.4375 59.8950 242.7075 60.4800 ;
		LAYER M3 ;
        RECT 242.4375 58.4400 242.7075 58.4700 ;
		LAYER M1 ;
        RECT 242.4375 59.4000 242.7075 59.4900 ;
		LAYER M3 ;
        RECT 242.4375 59.4300 242.7075 59.4600 ;
		LAYER M1 ;
        RECT 242.4375 58.9050 242.7075 58.9950 ;
		LAYER M2 ;
        RECT 242.4375 58.9350 242.7075 58.9650 ;
		LAYER VIA3 ;
        RECT 242.4375 59.4300 242.7075 59.4600 ;
		LAYER M2 ;
        RECT 242.4375 59.4300 242.7075 59.4600 ;
		LAYER M1 ;
        RECT 242.4375 119.4225 242.7075 119.5425 ;
		LAYER M3 ;
        RECT 242.4375 125.9175 242.7075 125.9475 ;
		LAYER M2 ;
        RECT 242.4375 125.9175 242.7075 125.9475 ;
		LAYER VIA3 ;
        RECT 242.4375 125.9175 242.7075 125.9475 ;
		LAYER VIA3 ;
        RECT 242.4375 119.4525 242.7075 119.5125 ;
		LAYER M1 ;
        RECT 242.4375 124.9200 242.7075 125.4825 ;
		LAYER M1 ;
        RECT 242.4375 118.9275 242.7075 119.0175 ;
		LAYER M3 ;
        RECT 242.4375 129.3975 242.7075 129.4275 ;
		LAYER M2 ;
        RECT 242.4375 129.3975 242.7075 129.4275 ;
		LAYER VIA3 ;
        RECT 242.4375 129.3975 242.7075 129.4275 ;
		LAYER M3 ;
        RECT 242.4375 118.9575 242.7075 118.9875 ;
		LAYER M1 ;
        RECT 242.4375 129.3675 242.7075 129.4575 ;
		LAYER VIA3 ;
        RECT 242.4375 129.8925 242.7075 129.9525 ;
		LAYER M3 ;
        RECT 242.4375 126.4125 242.7075 126.4725 ;
		LAYER VIA3 ;
        RECT 242.4375 126.4125 242.7075 126.4725 ;
		LAYER M3 ;
        RECT 242.4375 127.4325 242.7075 127.9650 ;
		LAYER M1 ;
        RECT 242.4375 126.3825 242.7075 126.5025 ;
		LAYER VIA3 ;
        RECT 242.4375 126.9375 242.7075 126.9675 ;
		LAYER M2 ;
        RECT 242.4375 127.4325 242.7075 127.9650 ;
		LAYER VIA3 ;
        RECT 242.4375 127.4325 242.7075 127.9650 ;
		LAYER M2 ;
        RECT 242.4375 126.4125 242.7075 126.4725 ;
		LAYER M1 ;
        RECT 242.4375 128.4000 242.7075 128.9625 ;
		LAYER M3 ;
        RECT 242.4375 128.4300 242.7075 128.9325 ;
		LAYER VIA3 ;
        RECT 242.4375 128.4300 242.7075 128.9325 ;
		LAYER VIA3 ;
        RECT 242.4375 130.4175 242.7075 130.4475 ;
		LAYER M3 ;
        RECT 242.4375 130.4175 242.7075 130.4475 ;
		LAYER M2 ;
        RECT 242.4375 129.8925 242.7075 129.9525 ;
		LAYER M3 ;
        RECT 242.4375 129.8925 242.7075 129.9525 ;
		LAYER M1 ;
        RECT 242.4375 129.8625 242.7075 129.9825 ;
		LAYER VIA3 ;
        RECT 242.4375 55.4400 242.7075 55.9425 ;
		LAYER M2 ;
        RECT 242.4375 55.4400 242.7075 55.9425 ;
		LAYER M1 ;
        RECT 242.4375 55.4100 242.7075 55.9725 ;
		LAYER M3 ;
        RECT 242.4375 54.4425 242.7075 54.9750 ;
		LAYER M2 ;
        RECT 242.4375 56.4075 242.7075 56.4375 ;
		LAYER M1 ;
        RECT 242.4375 56.3775 242.7075 56.4675 ;
		LAYER M1 ;
        RECT 242.4375 56.8725 242.7075 58.0050 ;
		LAYER M3 ;
        RECT 242.4375 56.4075 242.7075 56.4375 ;
		LAYER VIA3 ;
        RECT 242.4375 56.4075 242.7075 56.4375 ;
		LAYER VIA3 ;
        RECT 242.4375 50.9625 242.7075 51.4950 ;
		LAYER M2 ;
        RECT 242.4375 50.9625 242.7075 51.4950 ;
		LAYER M3 ;
        RECT 242.4375 50.9625 242.7075 51.4950 ;
		LAYER M1 ;
        RECT 242.4375 50.9325 242.7075 51.5250 ;
		LAYER M2 ;
        RECT 242.4375 50.4675 242.7075 50.4975 ;
		LAYER M3 ;
        RECT 242.4375 52.9275 242.7075 52.9575 ;
		LAYER M1 ;
        RECT 242.4375 52.8975 242.7075 52.9875 ;
		LAYER VIA3 ;
        RECT 242.4375 53.4225 242.7075 53.4825 ;
		LAYER M1 ;
        RECT 242.4375 53.3925 242.7075 53.5125 ;
		LAYER M1 ;
        RECT 242.4375 50.4375 242.7075 50.5275 ;
		LAYER VIA3 ;
        RECT 242.4375 50.4675 242.7075 50.4975 ;
		LAYER M3 ;
        RECT 242.4375 50.4675 242.7075 50.4975 ;
		LAYER M2 ;
        RECT 242.4375 51.9600 242.7075 52.4625 ;
		LAYER M3 ;
        RECT 242.4375 51.9600 242.7075 52.4625 ;
		LAYER VIA3 ;
        RECT 242.4375 51.9600 242.7075 52.4625 ;
		LAYER M1 ;
        RECT 242.4375 51.9300 242.7075 52.4925 ;
		LAYER M3 ;
        RECT 242.4375 137.3775 242.7075 137.4075 ;
		LAYER M2 ;
        RECT 242.4375 135.3900 242.7075 135.8925 ;
		LAYER M1 ;
        RECT 242.4375 136.3275 242.7075 136.4175 ;
		LAYER M3 ;
        RECT 242.4375 135.3900 242.7075 135.8925 ;
		LAYER VIA3 ;
        RECT 242.4375 135.3900 242.7075 135.8925 ;
		LAYER M2 ;
        RECT 242.4375 136.8525 242.7075 136.9125 ;
		LAYER M1 ;
        RECT 242.4375 136.8225 242.7075 136.9425 ;
		LAYER M2 ;
        RECT 242.4375 136.3575 242.7075 136.3875 ;
		LAYER M3 ;
        RECT 242.4375 136.3575 242.7075 136.3875 ;
		LAYER M2 ;
        RECT 242.4375 126.9375 242.7075 126.9675 ;
		LAYER VIA3 ;
        RECT 242.4375 0.0000 242.7075 1.2825 ;
		LAYER M2 ;
        RECT 242.4375 0.0000 242.7075 1.2825 ;
		LAYER M1 ;
        RECT 242.4375 1.7175 242.7075 1.8075 ;
		LAYER M4 ;
        RECT 242.2050 0.0000 242.7075 141.6150 ;
		LAYER M1 ;
        RECT 242.4375 2.2125 242.7075 2.8050 ;
		LAYER M1 ;
        RECT 242.4375 0.0000 242.7075 1.3125 ;
		LAYER M3 ;
        RECT 242.4375 0.0000 242.7075 1.2825 ;
		LAYER M1 ;
        RECT 242.4375 132.8475 242.7075 132.9375 ;
		LAYER M3 ;
        RECT 242.4375 138.8700 242.7075 139.3725 ;
		LAYER VIA3 ;
        RECT 242.4375 138.8700 242.7075 139.3725 ;
		LAYER VIA3 ;
        RECT 242.4375 137.3775 242.7075 137.4075 ;
		LAYER M3 ;
        RECT 242.4375 134.3925 242.7075 134.9250 ;
		LAYER M1 ;
        RECT 242.4375 135.3600 242.7075 135.9225 ;
		LAYER VIA3 ;
        RECT 242.4375 134.3925 242.7075 134.9250 ;
		LAYER M3 ;
        RECT 242.4375 136.8525 242.7075 136.9125 ;
		LAYER M3 ;
        RECT 242.4375 63.7500 242.7075 63.9750 ;
		LAYER M2 ;
        RECT 242.4375 139.8375 242.7075 139.8675 ;
		LAYER VIA3 ;
        RECT 242.4375 139.8375 242.7075 139.8675 ;
		LAYER M3 ;
        RECT 242.4375 1.7475 242.7075 1.7775 ;
		LAYER VIA3 ;
        RECT 242.4375 1.7475 242.7075 1.7775 ;
		LAYER M3 ;
        RECT 242.4375 62.1000 242.7075 62.3250 ;
		LAYER M3 ;
        RECT 242.4375 137.8725 242.7075 138.4050 ;
		LAYER M2 ;
        RECT 242.4375 137.8725 242.7075 138.4050 ;
		LAYER VIA3 ;
        RECT 242.4375 137.8725 242.7075 138.4050 ;
		LAYER M1 ;
        RECT 242.4375 137.8425 242.7075 138.4350 ;
	END
END SRAM2048x32M4_1001


MACRO TAPCELL_0010
    CLASS CORE ;
    FOREIGN TAPCELL_0010 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.0500 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.5025 -0.0750 1.0500 0.0750 ;
        RECT 0.3825 -0.0750 0.5025 0.3450 ;
        RECT 0.0000 -0.0750 0.3825 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.6525 0.9750 1.0500 1.1250 ;
        RECT 0.5325 0.5925 0.6525 1.1250 ;
        RECT 0.0000 0.9750 0.5325 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 0.5625 0.6225 0.6225 0.6825 ;
        RECT 0.5625 0.7875 0.6225 0.8475 ;
        RECT 0.4125 0.2550 0.4725 0.3150 ;
    END
END TAPCELL_0010


MACRO TIEH_0010
    CLASS CORE ;
    FOREIGN TIEH_0010 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.4200 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.3075 0.3675 0.3825 0.8325 ;
        RECT 0.2775 0.6675 0.3075 0.8325 ;
        END
    END Z
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.3675 -0.0750 0.4200 0.0750 ;
        RECT 0.2625 -0.0750 0.3675 0.2625 ;
        RECT 0.0000 -0.0750 0.2625 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.1425 0.9750 0.4200 1.1250 ;
        RECT 0.0675 0.8025 0.1425 1.1250 ;
        RECT 0.0000 0.9750 0.0675 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 0.2850 0.1800 0.3450 0.2400 ;
        RECT 0.2850 0.7200 0.3450 0.7800 ;
        RECT 0.1725 0.4800 0.2325 0.5400 ;
        RECT 0.0750 0.2175 0.1350 0.2775 ;
        RECT 0.0750 0.8325 0.1350 0.8925 ;
        LAYER M1 ;
        RECT 0.1425 0.4500 0.2325 0.5700 ;
        RECT 0.0675 0.1800 0.1425 0.5700 ;
    END
END TIEH_0010


MACRO TIEL_0010
    CLASS CORE ;
    FOREIGN TIEL_0010 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.4200 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.3075 0.2175 0.3825 0.6825 ;
        RECT 0.2775 0.2175 0.3075 0.3825 ;
        END
    END ZN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.1425 -0.0750 0.4200 0.0750 ;
        RECT 0.0675 -0.0750 0.1425 0.3000 ;
        RECT 0.0000 -0.0750 0.0675 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 0.3525 0.9750 0.4200 1.1250 ;
        RECT 0.2775 0.8025 0.3525 1.1250 ;
        RECT 0.0000 0.9750 0.2775 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 0.2850 0.2700 0.3450 0.3300 ;
        RECT 0.2850 0.8325 0.3450 0.8925 ;
        RECT 0.1725 0.4800 0.2325 0.5400 ;
        RECT 0.0750 0.2100 0.1350 0.2700 ;
        RECT 0.0750 0.7125 0.1350 0.7725 ;
        LAYER M1 ;
        RECT 0.1425 0.4500 0.2325 0.5700 ;
        RECT 0.0675 0.4500 0.1425 0.8175 ;
    END
END TIEL_0010


MACRO XNR2_0011
    CLASS CORE ;
    FOREIGN XNR2_0011 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.8900 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 1.7775 0.3075 1.8525 0.7350 ;
        RECT 1.6125 0.3075 1.7775 0.3825 ;
        RECT 1.6125 0.6600 1.7775 0.7350 ;
        RECT 1.5375 0.2175 1.6125 0.3825 ;
        RECT 1.5375 0.6600 1.6125 0.8325 ;
        END
    END ZN
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.2825 0.1125 1.7475 0.1875 ;
        RECT 1.1775 0.1125 1.2825 0.4800 ;
        VIA 1.2300 0.4050 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.4575 0.4950 0.9000 0.5700 ;
        RECT 0.2775 0.4950 0.4575 0.7875 ;
        RECT 0.1875 0.4950 0.2775 0.6150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.8450 -0.0750 1.8900 0.0750 ;
        RECT 1.7250 -0.0750 1.8450 0.2325 ;
        RECT 1.4025 -0.0750 1.7250 0.0750 ;
        RECT 1.3275 -0.0750 1.4025 0.2250 ;
        RECT 0.3750 -0.0750 1.3275 0.0750 ;
        RECT 0.2550 -0.0750 0.3750 0.2400 ;
        RECT 0.0000 -0.0750 0.2550 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.8450 0.9750 1.8900 1.1250 ;
        RECT 1.7250 0.8100 1.8450 1.1250 ;
        RECT 1.4175 0.9750 1.7250 1.1250 ;
        RECT 1.3125 0.7875 1.4175 1.1250 ;
        RECT 0.3750 0.9750 1.3125 1.1250 ;
        RECT 0.2550 0.8625 0.3750 1.1250 ;
        RECT 0.0000 0.9750 0.2550 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.7550 0.1725 1.8150 0.2325 ;
        RECT 1.7550 0.8175 1.8150 0.8775 ;
        RECT 1.6425 0.4875 1.7025 0.5475 ;
        RECT 1.5450 0.2700 1.6050 0.3300 ;
        RECT 1.5450 0.7200 1.6050 0.7800 ;
        RECT 1.4400 0.4875 1.5000 0.5475 ;
        RECT 1.3350 0.1350 1.3950 0.1950 ;
        RECT 1.3350 0.8175 1.3950 0.8775 ;
        RECT 1.2300 0.4575 1.2900 0.5175 ;
        RECT 1.1250 0.1800 1.1850 0.2400 ;
        RECT 1.1250 0.6675 1.1850 0.7275 ;
        RECT 1.0200 0.3750 1.0800 0.4350 ;
        RECT 0.9150 0.1725 0.9750 0.2325 ;
        RECT 0.9150 0.8250 0.9750 0.8850 ;
        RECT 0.6000 0.6600 0.6600 0.7200 ;
        RECT 0.3900 0.3450 0.4500 0.4050 ;
        RECT 0.3900 0.6600 0.4500 0.7200 ;
        RECT 0.2850 0.1650 0.3450 0.2250 ;
        RECT 0.2850 0.8700 0.3450 0.9300 ;
        RECT 0.1875 0.5250 0.2475 0.5850 ;
        RECT 0.0750 0.1875 0.1350 0.2475 ;
        RECT 0.0750 0.8175 0.1350 0.8775 ;
        RECT 0.8100 0.5025 0.8700 0.5625 ;
        RECT 0.7050 0.1725 0.7650 0.2325 ;
        RECT 0.7050 0.8325 0.7650 0.8925 ;
        LAYER M1 ;
        RECT 1.4625 0.4575 1.7025 0.5775 ;
        RECT 1.3725 0.4575 1.4625 0.6825 ;
        RECT 1.1625 0.3300 1.2975 0.5700 ;
        RECT 0.8625 0.1500 1.2150 0.2550 ;
        RECT 0.5625 0.6600 1.2150 0.7350 ;
        RECT 1.0050 0.3375 1.0875 0.4650 ;
        RECT 0.6225 0.8100 1.0200 0.9000 ;
        RECT 0.1575 0.3375 1.0050 0.4125 ;
        RECT 0.4650 0.1500 0.7875 0.2550 ;
        RECT 0.1125 0.7950 0.1650 0.9000 ;
        RECT 0.1125 0.1650 0.1575 0.4125 ;
        RECT 0.0525 0.1650 0.1125 0.9000 ;
        RECT 0.0375 0.3375 0.0525 0.9000 ;
        LAYER VIA1 ;
        RECT 1.3800 0.5625 1.4550 0.6375 ;
        RECT 0.9750 0.1650 1.0500 0.2400 ;
        RECT 0.9525 0.6600 1.0275 0.7350 ;
        RECT 0.7575 0.8100 0.8325 0.8850 ;
        RECT 0.6750 0.1650 0.7500 0.2400 ;
        LAYER M2 ;
        RECT 1.3575 0.5625 1.5300 0.6375 ;
        RECT 1.2825 0.5625 1.3575 0.9375 ;
        RECT 0.8325 0.8625 1.2825 0.9375 ;
        RECT 1.0125 0.1500 1.0875 0.2550 ;
        RECT 1.0125 0.6225 1.0425 0.7725 ;
        RECT 0.9375 0.1500 1.0125 0.7725 ;
        RECT 0.7575 0.1500 0.8325 0.9375 ;
        RECT 0.6375 0.1500 0.7575 0.2550 ;
    END
END XNR2_0011


MACRO XNR2_0111
    CLASS CORE ;
    FOREIGN XNR2_0111 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.3600 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 2.6775 0.2625 2.9925 0.7500 ;
        VIA 2.8350 0.3225 VIA12_slot ;
        VIA 2.8350 0.6675 VIA12_slot ;
        END
    END ZN
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 2.1675 0.2625 2.2425 0.6075 ;
        RECT 1.7025 0.2625 2.1675 0.3375 ;
        VIA 2.2050 0.5250 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.3125 0.3150 1.4175 0.5625 ;
        RECT 1.1175 0.3150 1.3125 0.3975 ;
        RECT 1.0350 0.2625 1.1175 0.3975 ;
        RECT 0.3975 0.2625 1.0350 0.3375 ;
        VIA 1.3650 0.4875 VIA12_square ;
        VIA 0.5100 0.3000 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 3.2925 -0.0750 3.3600 0.0750 ;
        RECT 3.2175 -0.0750 3.2925 0.3150 ;
        RECT 2.8950 -0.0750 3.2175 0.0750 ;
        RECT 2.7750 -0.0750 2.8950 0.1950 ;
        RECT 2.4525 -0.0750 2.7750 0.0750 ;
        RECT 2.3775 -0.0750 2.4525 0.3075 ;
        RECT 2.0625 -0.0750 2.3775 0.0750 ;
        RECT 1.9575 -0.0750 2.0625 0.2475 ;
        RECT 1.0050 -0.0750 1.9575 0.0750 ;
        RECT 0.8850 -0.0750 1.0050 0.1950 ;
        RECT 0.3525 -0.0750 0.8850 0.0750 ;
        RECT 0.2775 -0.0750 0.3525 0.3000 ;
        RECT 0.0000 -0.0750 0.2775 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 3.2925 0.9750 3.3600 1.1250 ;
        RECT 3.2175 0.6375 3.2925 1.1250 ;
        RECT 2.8875 0.9750 3.2175 1.1250 ;
        RECT 2.7825 0.8025 2.8875 1.1250 ;
        RECT 2.4750 0.9750 2.7825 1.1250 ;
        RECT 2.3550 0.6600 2.4750 1.1250 ;
        RECT 2.0550 0.9750 2.3550 1.1250 ;
        RECT 1.9350 0.8025 2.0550 1.1250 ;
        RECT 0.7875 0.9750 1.9350 1.1250 ;
        RECT 0.6825 0.8100 0.7875 1.1250 ;
        RECT 0.3600 0.9750 0.6825 1.1250 ;
        RECT 0.2550 0.8100 0.3600 1.1250 ;
        RECT 0.0000 0.9750 0.2550 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 3.2250 0.2250 3.2850 0.2850 ;
        RECT 3.2250 0.6675 3.2850 0.7275 ;
        RECT 3.2250 0.8325 3.2850 0.8925 ;
        RECT 3.1200 0.4650 3.1800 0.5250 ;
        RECT 3.0150 0.2250 3.0750 0.2850 ;
        RECT 3.0150 0.7575 3.0750 0.8175 ;
        RECT 2.9100 0.4650 2.9700 0.5250 ;
        RECT 2.8050 0.1275 2.8650 0.1875 ;
        RECT 2.8050 0.8325 2.8650 0.8925 ;
        RECT 2.7000 0.4650 2.7600 0.5250 ;
        RECT 2.5950 0.2250 2.6550 0.2850 ;
        RECT 2.5950 0.7575 2.6550 0.8175 ;
        RECT 2.4900 0.4650 2.5500 0.5250 ;
        RECT 2.3850 0.2175 2.4450 0.2775 ;
        RECT 2.3850 0.6675 2.4450 0.7275 ;
        RECT 2.3850 0.8325 2.4450 0.8925 ;
        RECT 2.2800 0.4875 2.3400 0.5475 ;
        RECT 2.1750 0.3075 2.2350 0.3675 ;
        RECT 2.1750 0.7275 2.2350 0.7875 ;
        RECT 2.0700 0.4875 2.1300 0.5475 ;
        RECT 1.9650 0.1575 2.0250 0.2175 ;
        RECT 1.9650 0.8100 2.0250 0.8700 ;
        RECT 1.7550 0.6525 1.8150 0.7125 ;
        RECT 1.6500 0.4500 1.7100 0.5100 ;
        RECT 1.5450 0.1725 1.6050 0.2325 ;
        RECT 1.5450 0.8250 1.6050 0.8850 ;
        RECT 1.4400 0.4800 1.5000 0.5400 ;
        RECT 1.3350 0.2325 1.3950 0.2925 ;
        RECT 1.3350 0.8175 1.3950 0.8775 ;
        RECT 1.2300 0.6450 1.2900 0.7050 ;
        RECT 1.1250 0.2400 1.1850 0.3000 ;
        RECT 1.1250 0.8175 1.1850 0.8775 ;
        RECT 1.0200 0.4950 1.0800 0.5550 ;
        RECT 0.9150 0.1275 0.9750 0.1875 ;
        RECT 0.8100 0.4950 0.8700 0.5550 ;
        RECT 0.7050 0.2775 0.7650 0.3375 ;
        RECT 0.7050 0.8325 0.7650 0.8925 ;
        RECT 0.6000 0.4800 0.6600 0.5400 ;
        RECT 0.4950 0.8250 0.5550 0.8850 ;
        RECT 0.3900 0.4800 0.4500 0.5400 ;
        RECT 0.2850 0.2025 0.3450 0.2625 ;
        RECT 0.2850 0.8400 0.3450 0.9000 ;
        RECT 0.1875 0.4650 0.2475 0.5250 ;
        RECT 0.0750 0.2325 0.1350 0.2925 ;
        RECT 0.0750 0.7350 0.1350 0.7950 ;
        LAYER M1 ;
        RECT 2.4375 0.4425 3.2100 0.5475 ;
        RECT 2.9925 0.1950 3.0975 0.3675 ;
        RECT 3.0075 0.6225 3.0825 0.8700 ;
        RECT 2.6625 0.6225 3.0075 0.7125 ;
        RECT 2.6775 0.2775 2.9925 0.3675 ;
        RECT 2.5725 0.1950 2.6775 0.3675 ;
        RECT 2.5875 0.6225 2.6625 0.8700 ;
        RECT 2.2575 0.4650 2.3625 0.5700 ;
        RECT 2.1900 0.2775 2.2650 0.3900 ;
        RECT 1.9950 0.4800 2.2575 0.5700 ;
        RECT 2.1675 0.6450 2.2425 0.8250 ;
        RECT 2.1450 0.2775 2.1900 0.3975 ;
        RECT 1.8825 0.6450 2.1675 0.7200 ;
        RECT 1.8825 0.3225 2.1450 0.3975 ;
        RECT 1.8075 0.1500 1.8825 0.7200 ;
        RECT 1.5225 0.1500 1.8075 0.2550 ;
        RECT 1.1925 0.6450 1.8075 0.7200 ;
        RECT 1.5975 0.3300 1.7325 0.5700 ;
        RECT 1.3125 0.7950 1.6575 0.9000 ;
        RECT 1.2450 0.4350 1.5225 0.5625 ;
        RECT 1.2675 0.1500 1.4250 0.3600 ;
        RECT 1.0875 0.7950 1.2075 0.9000 ;
        RECT 1.1175 0.1950 1.1925 0.3450 ;
        RECT 0.6525 0.2700 1.1175 0.3450 ;
        RECT 0.7950 0.4650 1.0950 0.5850 ;
        RECT 1.0125 0.6600 1.0875 0.9000 ;
        RECT 0.6075 0.6600 1.0125 0.7350 ;
        RECT 0.5475 0.4500 0.6900 0.5550 ;
        RECT 0.5325 0.6600 0.6075 0.9000 ;
        RECT 0.4725 0.2175 0.5475 0.5550 ;
        RECT 0.4650 0.8100 0.5325 0.9000 ;
        RECT 0.1875 0.4350 0.4725 0.5550 ;
        RECT 0.1500 0.6300 0.4575 0.7350 ;
        RECT 0.1125 0.6300 0.1500 0.8325 ;
        RECT 0.1125 0.2025 0.1425 0.3225 ;
        RECT 0.0375 0.2025 0.1125 0.8325 ;
        LAYER VIA1 ;
        RECT 2.4825 0.4575 2.5575 0.5325 ;
        RECT 1.6275 0.4125 1.7025 0.4875 ;
        RECT 1.4625 0.8100 1.5375 0.8850 ;
        RECT 1.3125 0.1650 1.3875 0.2400 ;
        RECT 0.9075 0.5100 0.9825 0.5850 ;
        RECT 0.3450 0.6450 0.4200 0.7200 ;
        LAYER M2 ;
        RECT 2.4375 0.4200 2.5725 0.5700 ;
        RECT 2.3625 0.1125 2.4375 0.8850 ;
        RECT 1.5375 0.1125 2.3625 0.1875 ;
        RECT 1.4175 0.8100 2.3625 0.8850 ;
        RECT 1.6125 0.4125 1.7775 0.4875 ;
        RECT 1.5375 0.4125 1.6125 0.7200 ;
        RECT 1.4550 0.1125 1.5375 0.2400 ;
        RECT 0.9975 0.6450 1.5375 0.7200 ;
        RECT 1.2675 0.1650 1.4550 0.2400 ;
        RECT 0.8925 0.4725 0.9975 0.7200 ;
        RECT 0.2700 0.6450 0.8925 0.7200 ;
    END
END XNR2_0111


MACRO XNR2_1000
    CLASS CORE ;
    FOREIGN XNR2_1000 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.5100 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 5.8800 0.3150 6.0375 0.4350 ;
        RECT 5.8800 0.6150 6.0375 0.7350 ;
        RECT 5.5650 0.3150 5.8800 0.7350 ;
        RECT 5.4075 0.3150 5.5650 0.4350 ;
        RECT 5.4075 0.6150 5.5650 0.7350 ;
        VIA 5.8800 0.3750 VIA12_slot ;
        VIA 5.8800 0.6750 VIA12_slot ;
        VIA 5.5650 0.3750 VIA12_slot ;
        VIA 5.5650 0.6750 VIA12_slot ;
        END
    END ZN
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.1100 0.4350 1.2225 0.6375 ;
        RECT 0.6000 0.5625 1.1100 0.6375 ;
        VIA 1.1700 0.5175 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 3.2325 0.4125 3.9975 0.4875 ;
        RECT 3.1275 0.4125 3.2325 0.6075 ;
        VIA 3.8775 0.4500 VIA12_square ;
        VIA 3.1800 0.5175 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 3.5400 -0.0750 6.5100 0.0750 ;
        RECT 3.3900 -0.0750 3.5400 0.2175 ;
        RECT 3.1050 -0.0750 3.3900 0.0750 ;
        RECT 2.9850 -0.0750 3.1050 0.2250 ;
        RECT 2.6850 -0.0750 2.9850 0.0750 ;
        RECT 2.5650 -0.0750 2.6850 0.2325 ;
        RECT 2.2650 -0.0750 2.5650 0.0750 ;
        RECT 2.1450 -0.0750 2.2650 0.2325 ;
        RECT 1.8450 -0.0750 2.1450 0.0750 ;
        RECT 1.7250 -0.0750 1.8450 0.2325 ;
        RECT 1.4250 -0.0750 1.7250 0.0750 ;
        RECT 1.3050 -0.0750 1.4250 0.2325 ;
        RECT 1.0050 -0.0750 1.3050 0.0750 ;
        RECT 0.8850 -0.0750 1.0050 0.2325 ;
        RECT 0.5775 -0.0750 0.8850 0.0750 ;
        RECT 0.4725 -0.0750 0.5775 0.2325 ;
        RECT 0.1650 -0.0750 0.4725 0.0750 ;
        RECT 0.0450 -0.0750 0.1650 0.2325 ;
        RECT 0.0000 -0.0750 0.0450 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 3.5250 0.9750 6.5100 1.1250 ;
        RECT 3.4050 0.8325 3.5250 1.1250 ;
        RECT 3.1200 0.9750 3.4050 1.1250 ;
        RECT 2.9700 0.8325 3.1200 1.1250 ;
        RECT 2.6850 0.9750 2.9700 1.1250 ;
        RECT 2.5650 0.8400 2.6850 1.1250 ;
        RECT 2.2650 0.9750 2.5650 1.1250 ;
        RECT 2.1450 0.8400 2.2650 1.1250 ;
        RECT 1.8450 0.9750 2.1450 1.1250 ;
        RECT 1.7250 0.8400 1.8450 1.1250 ;
        RECT 1.4250 0.9750 1.7250 1.1250 ;
        RECT 1.3050 0.8400 1.4250 1.1250 ;
        RECT 1.0050 0.9750 1.3050 1.1250 ;
        RECT 0.8850 0.8400 1.0050 1.1250 ;
        RECT 0.5850 0.9750 0.8850 1.1250 ;
        RECT 0.4650 0.8400 0.5850 1.1250 ;
        RECT 0.1650 0.9750 0.4650 1.1250 ;
        RECT 0.0450 0.8100 0.1650 1.1250 ;
        RECT 0.0000 0.9750 0.0450 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 6.3750 0.3075 6.4350 0.3675 ;
        RECT 6.3750 0.6750 6.4350 0.7350 ;
        RECT 6.2700 0.4950 6.3300 0.5550 ;
        RECT 6.1650 0.1575 6.2250 0.2175 ;
        RECT 6.1650 0.8325 6.2250 0.8925 ;
        RECT 6.0600 0.4950 6.1200 0.5550 ;
        RECT 5.9550 0.3225 6.0150 0.3825 ;
        RECT 5.9550 0.6750 6.0150 0.7350 ;
        RECT 5.8500 0.4950 5.9100 0.5550 ;
        RECT 5.7450 0.1575 5.8050 0.2175 ;
        RECT 5.7450 0.8325 5.8050 0.8925 ;
        RECT 5.6400 0.4950 5.7000 0.5550 ;
        RECT 5.5350 0.3225 5.5950 0.3825 ;
        RECT 5.5350 0.6750 5.5950 0.7350 ;
        RECT 5.4300 0.4950 5.4900 0.5550 ;
        RECT 5.3250 0.1575 5.3850 0.2175 ;
        RECT 5.3250 0.8325 5.3850 0.8925 ;
        RECT 5.2200 0.4950 5.2800 0.5550 ;
        RECT 5.1150 0.2625 5.1750 0.3225 ;
        RECT 5.1150 0.6750 5.1750 0.7350 ;
        RECT 5.0100 0.4800 5.0700 0.5400 ;
        RECT 4.9050 0.3000 4.9650 0.3600 ;
        RECT 4.9050 0.6675 4.9650 0.7275 ;
        RECT 4.8000 0.4800 4.8600 0.5400 ;
        RECT 4.6950 0.1575 4.7550 0.2175 ;
        RECT 4.6950 0.8325 4.7550 0.8925 ;
        RECT 4.5900 0.4800 4.6500 0.5400 ;
        RECT 4.4850 0.3000 4.5450 0.3600 ;
        RECT 4.4850 0.6675 4.5450 0.7275 ;
        RECT 4.3800 0.4800 4.4400 0.5400 ;
        RECT 4.2750 0.1575 4.3350 0.2175 ;
        RECT 4.2750 0.8325 4.3350 0.8925 ;
        RECT 4.1700 0.4800 4.2300 0.5400 ;
        RECT 4.0650 0.3000 4.1250 0.3600 ;
        RECT 4.0650 0.6825 4.1250 0.7425 ;
        RECT 3.9600 0.4800 4.0200 0.5400 ;
        RECT 3.8550 0.1875 3.9150 0.2475 ;
        RECT 3.8550 0.8025 3.9150 0.8625 ;
        RECT 3.6450 0.3075 3.7050 0.3675 ;
        RECT 3.6450 0.6900 3.7050 0.7500 ;
        RECT 3.5400 0.4875 3.6000 0.5475 ;
        RECT 3.4350 0.1575 3.4950 0.2175 ;
        RECT 3.4350 0.8325 3.4950 0.8925 ;
        RECT 3.3300 0.4875 3.3900 0.5475 ;
        RECT 3.2250 0.3075 3.2850 0.3675 ;
        RECT 3.2250 0.6900 3.2850 0.7500 ;
        RECT 3.1200 0.4875 3.1800 0.5475 ;
        RECT 3.0150 0.1425 3.0750 0.2025 ;
        RECT 3.0150 0.8325 3.0750 0.8925 ;
        RECT 2.9100 0.4875 2.9700 0.5475 ;
        RECT 2.8050 0.2925 2.8650 0.3525 ;
        RECT 2.8050 0.7200 2.8650 0.7800 ;
        RECT 2.7000 0.4875 2.7600 0.5475 ;
        RECT 2.5950 0.1650 2.6550 0.2250 ;
        RECT 2.5950 0.8475 2.6550 0.9075 ;
        RECT 2.4900 0.4875 2.5500 0.5475 ;
        RECT 2.3850 0.3075 2.4450 0.3675 ;
        RECT 2.3850 0.6900 2.4450 0.7500 ;
        RECT 2.2800 0.4875 2.3400 0.5475 ;
        RECT 2.1750 0.1650 2.2350 0.2250 ;
        RECT 2.1750 0.8475 2.2350 0.9075 ;
        RECT 2.0700 0.4875 2.1300 0.5475 ;
        RECT 1.9650 0.2925 2.0250 0.3525 ;
        RECT 1.9650 0.7350 2.0250 0.7950 ;
        RECT 1.8600 0.4875 1.9200 0.5475 ;
        RECT 1.7550 0.1650 1.8150 0.2250 ;
        RECT 1.7550 0.8475 1.8150 0.9075 ;
        RECT 1.6500 0.4875 1.7100 0.5475 ;
        RECT 1.5450 0.3075 1.6050 0.3675 ;
        RECT 1.5450 0.6900 1.6050 0.7500 ;
        RECT 1.4400 0.4875 1.5000 0.5475 ;
        RECT 1.3350 0.1650 1.3950 0.2250 ;
        RECT 1.3350 0.8475 1.3950 0.9075 ;
        RECT 1.2300 0.4875 1.2900 0.5475 ;
        RECT 1.1250 0.3075 1.1850 0.3675 ;
        RECT 1.1250 0.6900 1.1850 0.7500 ;
        RECT 1.0200 0.4875 1.0800 0.5475 ;
        RECT 0.9150 0.1650 0.9750 0.2250 ;
        RECT 0.9150 0.8475 0.9750 0.9075 ;
        RECT 0.8100 0.4875 0.8700 0.5475 ;
        RECT 0.7050 0.3075 0.7650 0.3675 ;
        RECT 0.7050 0.6900 0.7650 0.7500 ;
        RECT 0.6000 0.4875 0.6600 0.5475 ;
        RECT 0.4950 0.1500 0.5550 0.2100 ;
        RECT 0.4950 0.8475 0.5550 0.9075 ;
        RECT 0.3900 0.4875 0.4500 0.5475 ;
        RECT 0.2850 0.2925 0.3450 0.3525 ;
        RECT 0.2850 0.7350 0.3450 0.7950 ;
        RECT 0.1800 0.4875 0.2400 0.5475 ;
        RECT 0.0750 0.1650 0.1350 0.2250 ;
        RECT 0.0750 0.8175 0.1350 0.8775 ;
        LAYER M1 ;
        RECT 6.3450 0.2775 6.4650 0.4125 ;
        RECT 6.3600 0.6375 6.4425 0.7875 ;
        RECT 5.3400 0.4875 6.3900 0.5625 ;
        RECT 5.4075 0.6375 6.3600 0.7350 ;
        RECT 5.4075 0.3075 6.3450 0.4125 ;
        RECT 5.4525 0.1500 6.2775 0.2250 ;
        RECT 5.4075 0.8250 6.2550 0.9000 ;
        RECT 5.2875 0.1500 5.4525 0.2325 ;
        RECT 5.1825 0.3075 5.4075 0.3825 ;
        RECT 5.1375 0.6600 5.4075 0.7350 ;
        RECT 5.2425 0.8175 5.4075 0.9000 ;
        RECT 5.1450 0.4575 5.3400 0.5850 ;
        RECT 5.1075 0.1500 5.1825 0.3825 ;
        RECT 5.0625 0.6600 5.1375 0.9000 ;
        RECT 3.9300 0.1500 5.1075 0.2250 ;
        RECT 4.9650 0.4500 5.0700 0.5700 ;
        RECT 3.9225 0.8250 5.0625 0.9000 ;
        RECT 4.0350 0.3000 4.9950 0.3750 ;
        RECT 4.4025 0.6450 4.9875 0.7500 ;
        RECT 3.9300 0.4500 4.9650 0.5400 ;
        RECT 4.0350 0.6750 4.4025 0.7500 ;
        RECT 3.8250 0.1500 3.9300 0.2850 ;
        RECT 3.8250 0.3750 3.9300 0.5400 ;
        RECT 3.8475 0.7575 3.9225 0.9000 ;
        RECT 3.6750 0.3075 3.7500 0.7575 ;
        RECT 3.1875 0.3075 3.6750 0.3825 ;
        RECT 3.1875 0.6525 3.6750 0.7575 ;
        RECT 3.0825 0.4575 3.6000 0.5775 ;
        RECT 2.8725 0.3000 3.0750 0.3825 ;
        RECT 2.8425 0.4725 3.0000 0.5775 ;
        RECT 2.7975 0.2625 2.8725 0.3825 ;
        RECT 2.7975 0.6825 2.8725 0.8175 ;
        RECT 1.8600 0.4575 2.8425 0.5775 ;
        RECT 2.0325 0.3075 2.7975 0.3825 ;
        RECT 2.0325 0.6825 2.7975 0.7575 ;
        RECT 1.9575 0.2250 2.0325 0.3825 ;
        RECT 1.9575 0.6825 2.0325 0.8400 ;
        RECT 1.7850 0.3075 1.8600 0.7575 ;
        RECT 0.3525 0.3075 1.7850 0.3825 ;
        RECT 0.3525 0.6825 1.7850 0.7575 ;
        RECT 0.1500 0.4575 1.7100 0.5775 ;
        RECT 0.2775 0.2325 0.3525 0.3825 ;
        RECT 0.2775 0.6825 0.3525 0.8400 ;
        LAYER VIA1 ;
        RECT 5.3325 0.1575 5.4075 0.2325 ;
        RECT 5.2875 0.8175 5.3625 0.8925 ;
        RECT 5.1825 0.4800 5.2575 0.5550 ;
        RECT 4.4475 0.6675 4.5225 0.7425 ;
        RECT 4.2225 0.3000 4.2975 0.3750 ;
        RECT 3.6750 0.5625 3.7500 0.6375 ;
        RECT 2.9550 0.3075 3.0300 0.3825 ;
        RECT 2.7975 0.4875 2.8725 0.5625 ;
        RECT 2.5875 0.6825 2.6625 0.7575 ;
        RECT 2.5125 0.3075 2.5875 0.3825 ;
        LAYER M2 ;
        RECT 5.9100 0.3150 6.0375 0.4350 ;
        RECT 5.9100 0.6150 6.0375 0.7350 ;
        RECT 5.4075 0.3150 5.5350 0.4350 ;
        RECT 5.4075 0.6150 5.5350 0.7350 ;
        RECT 5.2875 0.1125 5.4525 0.2325 ;
        RECT 5.2425 0.8175 5.4075 0.9375 ;
        RECT 2.8725 0.1125 5.2875 0.1875 ;
        RECT 5.1825 0.4275 5.2575 0.6225 ;
        RECT 2.6625 0.8625 5.2425 0.9375 ;
        RECT 4.5375 0.4275 5.1825 0.5025 ;
        RECT 4.4325 0.6225 4.5450 0.7875 ;
        RECT 4.4625 0.4275 4.5375 0.5475 ;
        RECT 4.3575 0.4725 4.4625 0.5475 ;
        RECT 2.8725 0.7125 4.4325 0.7875 ;
        RECT 4.2825 0.4725 4.3575 0.6375 ;
        RECT 4.1775 0.2625 4.3425 0.3900 ;
        RECT 3.6150 0.5625 4.2825 0.6375 ;
        RECT 3.0300 0.2625 4.1775 0.3375 ;
        RECT 2.9550 0.2625 3.0300 0.4500 ;
        RECT 2.7975 0.1125 2.8725 0.7875 ;
        RECT 2.5875 0.3075 2.6625 0.9375 ;
        RECT 2.4375 0.3075 2.5875 0.3825 ;
    END
END XNR2_1000


MACRO XNR2_1010
    CLASS CORE ;
    FOREIGN XNR2_1010 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.4700 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 0.7800 0.8625 1.2450 0.9375 ;
        RECT 0.7050 0.1500 0.7800 0.9375 ;
        RECT 0.6300 0.1500 0.7050 0.2550 ;
        VIA 0.7425 0.8475 VIA12_square ;
        VIA 0.7050 0.2025 VIA12_square ;
        END
    END ZN
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.3125 0.3675 1.4175 0.6825 ;
        RECT 1.2300 0.3675 1.3125 0.5550 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.1200 0.4125 0.5850 0.4875 ;
        VIA 0.2925 0.4500 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.4025 -0.0750 1.4700 0.0750 ;
        RECT 1.2975 -0.0750 1.4025 0.2550 ;
        RECT 0.3750 -0.0750 1.2975 0.0750 ;
        RECT 0.2550 -0.0750 0.3750 0.1875 ;
        RECT 0.0000 -0.0750 0.2550 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.4250 0.9750 1.4700 1.1250 ;
        RECT 1.3050 0.7875 1.4250 1.1250 ;
        RECT 0.3750 0.9750 1.3050 1.1250 ;
        RECT 0.2550 0.8700 0.3750 1.1250 ;
        RECT 0.0000 0.9750 0.2550 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.3350 0.1650 1.3950 0.2250 ;
        RECT 1.3350 0.7875 1.3950 0.8475 ;
        RECT 1.2300 0.4650 1.2900 0.5250 ;
        RECT 1.1250 0.1800 1.1850 0.2400 ;
        RECT 1.1250 0.7275 1.1850 0.7875 ;
        RECT 1.0200 0.4650 1.0800 0.5250 ;
        RECT 0.9150 0.1800 0.9750 0.2400 ;
        RECT 0.9150 0.8325 0.9750 0.8925 ;
        RECT 0.8100 0.5025 0.8700 0.5625 ;
        RECT 0.7050 0.1800 0.7650 0.2400 ;
        RECT 0.7050 0.8325 0.7650 0.8925 ;
        RECT 0.6000 0.6525 0.6600 0.7125 ;
        RECT 0.3975 0.6600 0.4575 0.7200 ;
        RECT 0.3900 0.3450 0.4500 0.4050 ;
        RECT 0.2850 0.1200 0.3450 0.1800 ;
        RECT 0.2850 0.8700 0.3450 0.9300 ;
        RECT 0.1875 0.4800 0.2475 0.5400 ;
        RECT 0.0750 0.1800 0.1350 0.2400 ;
        RECT 0.0750 0.8175 0.1350 0.8775 ;
        LAYER M1 ;
        RECT 0.8700 0.1500 1.2225 0.2550 ;
        RECT 1.1100 0.6600 1.1850 0.8250 ;
        RECT 0.6825 0.6600 1.1100 0.7350 ;
        RECT 1.0125 0.3300 1.0875 0.5550 ;
        RECT 0.3450 0.3300 1.0125 0.4050 ;
        RECT 0.5775 0.8100 1.0050 0.9000 ;
        RECT 0.7725 0.4800 0.8925 0.5850 ;
        RECT 0.4725 0.1500 0.7950 0.2550 ;
        RECT 0.5025 0.4800 0.7725 0.5550 ;
        RECT 0.5775 0.6300 0.6825 0.7350 ;
        RECT 0.4275 0.4800 0.5025 0.7275 ;
        RECT 0.1575 0.6525 0.4275 0.7275 ;
        RECT 0.2325 0.3300 0.3450 0.5775 ;
        RECT 0.1875 0.4500 0.2325 0.5775 ;
        RECT 0.1125 0.6525 0.1575 0.9000 ;
        RECT 0.1125 0.1500 0.1425 0.2700 ;
        RECT 0.0375 0.1500 0.1125 0.9000 ;
        LAYER VIA1 ;
        RECT 0.9075 0.1650 0.9825 0.2400 ;
        RECT 0.9075 0.6600 0.9825 0.7350 ;
        LAYER M2 ;
        RECT 0.9675 0.1275 0.9975 0.2775 ;
        RECT 0.9675 0.6225 0.9975 0.7725 ;
        RECT 0.8925 0.1275 0.9675 0.7725 ;
    END
END XNR2_1010


MACRO XNR3_0011
    CLASS CORE ;
    FOREIGN XNR3_0011 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.3600 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 3.2475 0.3075 3.3225 0.7350 ;
        RECT 3.0825 0.3075 3.2475 0.3825 ;
        RECT 3.0825 0.6600 3.2475 0.7350 ;
        RECT 3.0075 0.2175 3.0825 0.3825 ;
        RECT 3.0075 0.6600 3.0825 0.8325 ;
        END
    END ZN
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 2.7750 0.1125 3.0900 0.1875 ;
        RECT 2.7000 0.1125 2.7750 0.4875 ;
        RECT 2.3850 0.4125 2.7000 0.4875 ;
        VIA 2.6850 0.4500 VIA12_square ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.2150 0.5625 1.6800 0.6375 ;
        VIA 1.3575 0.6000 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.6075 0.3375 0.7800 0.4425 ;
        RECT 0.5325 0.3375 0.6075 0.6375 ;
        RECT 0.0675 0.5625 0.5325 0.6375 ;
        VIA 0.6975 0.3750 VIA12_square ;
        VIA 0.2700 0.6000 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 3.3150 -0.0750 3.3600 0.0750 ;
        RECT 3.1950 -0.0750 3.3150 0.2325 ;
        RECT 2.8875 -0.0750 3.1950 0.0750 ;
        RECT 2.7825 -0.0750 2.8875 0.2550 ;
        RECT 1.8450 -0.0750 2.7825 0.0750 ;
        RECT 1.7250 -0.0750 1.8450 0.2400 ;
        RECT 1.4100 -0.0750 1.7250 0.0750 ;
        RECT 1.3200 -0.0750 1.4100 0.2625 ;
        RECT 0.3675 -0.0750 1.3200 0.0750 ;
        RECT 0.2625 -0.0750 0.3675 0.2475 ;
        RECT 0.0000 -0.0750 0.2625 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 3.3150 0.9750 3.3600 1.1250 ;
        RECT 3.1950 0.8100 3.3150 1.1250 ;
        RECT 2.8950 0.9750 3.1950 1.1250 ;
        RECT 2.7900 0.8100 2.8950 1.1250 ;
        RECT 1.8450 0.9750 2.7900 1.1250 ;
        RECT 1.7250 0.8250 1.8450 1.1250 ;
        RECT 1.4025 0.9750 1.7250 1.1250 ;
        RECT 1.3275 0.7875 1.4025 1.1250 ;
        RECT 0.3675 0.9750 1.3275 1.1250 ;
        RECT 0.2625 0.8250 0.3675 1.1250 ;
        RECT 0.0000 0.9750 0.2625 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 3.2250 0.1725 3.2850 0.2325 ;
        RECT 3.2250 0.8175 3.2850 0.8775 ;
        RECT 3.1125 0.4875 3.1725 0.5475 ;
        RECT 3.0150 0.2700 3.0750 0.3300 ;
        RECT 3.0150 0.7200 3.0750 0.7800 ;
        RECT 2.9100 0.4875 2.9700 0.5475 ;
        RECT 2.8050 0.1650 2.8650 0.2250 ;
        RECT 2.8050 0.8400 2.8650 0.9000 ;
        RECT 2.7000 0.4650 2.7600 0.5250 ;
        RECT 2.5950 0.1800 2.6550 0.2400 ;
        RECT 2.5950 0.6600 2.6550 0.7200 ;
        RECT 2.4900 0.4500 2.5500 0.5100 ;
        RECT 2.3850 0.1800 2.4450 0.2400 ;
        RECT 2.3850 0.8325 2.4450 0.8925 ;
        RECT 2.2800 0.5025 2.3400 0.5625 ;
        RECT 2.1750 0.1800 2.2350 0.2400 ;
        RECT 2.1750 0.8325 2.2350 0.8925 ;
        RECT 2.0700 0.6600 2.1300 0.7200 ;
        RECT 1.8600 0.3600 1.9200 0.4200 ;
        RECT 1.8600 0.6300 1.9200 0.6900 ;
        RECT 1.7550 0.1575 1.8150 0.2175 ;
        RECT 1.7550 0.8550 1.8150 0.9150 ;
        RECT 1.6500 0.5250 1.7100 0.5850 ;
        RECT 1.5450 0.1800 1.6050 0.2400 ;
        RECT 1.5450 0.7950 1.6050 0.8550 ;
        RECT 1.3350 0.1725 1.3950 0.2325 ;
        RECT 1.3350 0.8175 1.3950 0.8775 ;
        RECT 1.2300 0.5100 1.2900 0.5700 ;
        RECT 1.1250 0.1800 1.1850 0.2400 ;
        RECT 1.1250 0.7200 1.1850 0.7800 ;
        RECT 1.0200 0.4950 1.0800 0.5550 ;
        RECT 0.9150 0.1725 0.9750 0.2325 ;
        RECT 0.9150 0.8325 0.9750 0.8925 ;
        RECT 0.8100 0.3525 0.8700 0.4125 ;
        RECT 0.7050 0.1650 0.7650 0.2250 ;
        RECT 0.7050 0.8325 0.7650 0.8925 ;
        RECT 0.6000 0.6600 0.6600 0.7200 ;
        RECT 0.3900 0.4200 0.4500 0.4800 ;
        RECT 0.3900 0.6600 0.4500 0.7200 ;
        RECT 0.2850 0.1575 0.3450 0.2175 ;
        RECT 0.2850 0.8475 0.3450 0.9075 ;
        RECT 0.1875 0.5175 0.2475 0.5775 ;
        RECT 0.0750 0.2700 0.1350 0.3300 ;
        RECT 0.0750 0.8175 0.1350 0.8775 ;
        LAYER M1 ;
        RECT 2.9325 0.4575 3.1725 0.5775 ;
        RECT 2.8425 0.4575 2.9325 0.6825 ;
        RECT 2.6325 0.3300 2.7675 0.5700 ;
        RECT 2.4825 0.1500 2.6925 0.2550 ;
        RECT 2.5650 0.6450 2.6850 0.7500 ;
        RECT 2.0400 0.6450 2.5650 0.7350 ;
        RECT 2.4825 0.3450 2.5575 0.5400 ;
        RECT 2.3100 0.1500 2.4825 0.2700 ;
        RECT 1.6275 0.3450 2.4825 0.4200 ;
        RECT 2.1000 0.8100 2.4750 0.9000 ;
        RECT 1.9350 0.4950 2.3775 0.5700 ;
        RECT 1.9275 0.1500 2.2350 0.2700 ;
        RECT 1.8300 0.4950 1.9350 0.7200 ;
        RECT 1.6425 0.4950 1.8300 0.6150 ;
        RECT 1.5675 0.7725 1.6350 0.8775 ;
        RECT 1.5675 0.1500 1.6275 0.4200 ;
        RECT 1.5225 0.1500 1.5675 0.8775 ;
        RECT 1.4850 0.3450 1.5225 0.8775 ;
        RECT 1.3050 0.4875 1.4100 0.6825 ;
        RECT 1.1925 0.4875 1.3050 0.5925 ;
        RECT 1.0500 0.1500 1.2075 0.4125 ;
        RECT 1.1175 0.6675 1.1925 0.8100 ;
        RECT 0.6900 0.6675 1.1175 0.7425 ;
        RECT 1.0050 0.4875 1.1100 0.5925 ;
        RECT 0.8850 0.1500 1.0500 0.2550 ;
        RECT 0.4575 0.4875 1.0050 0.5625 ;
        RECT 0.5850 0.8175 1.0050 0.9000 ;
        RECT 0.5625 0.3300 0.9450 0.4125 ;
        RECT 0.4650 0.1500 0.7950 0.2550 ;
        RECT 0.5775 0.6375 0.6900 0.7425 ;
        RECT 0.3675 0.6375 0.4800 0.7425 ;
        RECT 0.3825 0.3375 0.4575 0.5625 ;
        RECT 0.1425 0.3375 0.3825 0.4125 ;
        RECT 0.3075 0.6375 0.3675 0.7200 ;
        RECT 0.2325 0.4875 0.3075 0.7200 ;
        RECT 0.1875 0.4875 0.2325 0.6075 ;
        RECT 0.1125 0.7950 0.1575 0.9000 ;
        RECT 0.1125 0.2400 0.1425 0.4125 ;
        RECT 0.0375 0.2400 0.1125 0.9000 ;
        LAYER VIA1 ;
        RECT 2.8425 0.5625 2.9175 0.6375 ;
        RECT 2.4075 0.6450 2.4825 0.7200 ;
        RECT 2.3475 0.1725 2.4225 0.2475 ;
        RECT 2.2575 0.8100 2.3325 0.8850 ;
        RECT 1.9875 0.1800 2.0625 0.2550 ;
        RECT 1.8375 0.4950 1.9125 0.5700 ;
        RECT 1.0875 0.3225 1.1625 0.3975 ;
        RECT 1.0200 0.6675 1.0950 0.7425 ;
        RECT 0.8250 0.8175 0.9000 0.8925 ;
        RECT 0.5100 0.1725 0.5850 0.2475 ;
        LAYER M2 ;
        RECT 2.8425 0.5625 2.9925 0.6375 ;
        RECT 2.7675 0.5625 2.8425 0.8850 ;
        RECT 2.1150 0.8100 2.7675 0.8850 ;
        RECT 2.2650 0.6450 2.5275 0.7200 ;
        RECT 2.2650 0.1725 2.4675 0.2475 ;
        RECT 2.1900 0.1725 2.2650 0.7200 ;
        RECT 2.0400 0.1650 2.1150 0.8850 ;
        RECT 1.9500 0.1650 2.0400 0.2700 ;
        RECT 1.8375 0.4125 1.9125 0.6450 ;
        RECT 1.4325 0.4125 1.8375 0.4875 ;
        RECT 1.3575 0.1575 1.4325 0.4875 ;
        RECT 0.9450 0.1575 1.3575 0.2325 ;
        RECT 1.0950 0.3150 1.2075 0.4200 ;
        RECT 1.0200 0.3150 1.0950 0.7950 ;
        RECT 0.8700 0.1575 0.9450 0.9000 ;
        RECT 0.6225 0.1575 0.8700 0.2325 ;
        RECT 0.7800 0.8100 0.8700 0.9000 ;
        RECT 0.4725 0.1575 0.6225 0.2625 ;
    END
END XNR3_0011


MACRO XNR3_0111
    CLASS CORE ;
    FOREIGN XNR3_0111 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.2000 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 3.5175 0.2625 3.8325 0.7275 ;
        VIA 3.6750 0.3225 VIA12_slot ;
        VIA 3.6750 0.6675 VIA12_slot ;
        END
    END ZN
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 3.3375 0.6825 3.4425 0.7875 ;
        RECT 2.9625 0.7125 3.3375 0.7875 ;
        VIA 3.2550 0.7500 VIA12_square ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.2150 0.5625 1.6800 0.6375 ;
        VIA 1.3275 0.6000 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.6900 0.3375 0.7800 0.4425 ;
        RECT 0.6150 0.3375 0.6900 0.6375 ;
        RECT 0.1575 0.5625 0.6150 0.6375 ;
        VIA 0.6975 0.3750 VIA12_square ;
        VIA 0.2700 0.6000 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 4.1475 -0.0750 4.2000 0.0750 ;
        RECT 4.0425 -0.0750 4.1475 0.3000 ;
        RECT 3.7350 -0.0750 4.0425 0.0750 ;
        RECT 3.6150 -0.0750 3.7350 0.1950 ;
        RECT 3.3150 -0.0750 3.6150 0.0750 ;
        RECT 3.2250 -0.0750 3.3150 0.2925 ;
        RECT 2.2650 -0.0750 3.2250 0.0750 ;
        RECT 2.1450 -0.0750 2.2650 0.1875 ;
        RECT 1.4025 -0.0750 2.1450 0.0750 ;
        RECT 1.3200 -0.0750 1.4025 0.3150 ;
        RECT 0.3675 -0.0750 1.3200 0.0750 ;
        RECT 0.2625 -0.0750 0.3675 0.2475 ;
        RECT 0.0000 -0.0750 0.2625 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 4.1550 0.9750 4.2000 1.1250 ;
        RECT 4.0350 0.7725 4.1550 1.1250 ;
        RECT 3.7350 0.9750 4.0350 1.1250 ;
        RECT 3.6150 0.8175 3.7350 1.1250 ;
        RECT 3.3150 0.9750 3.6150 1.1250 ;
        RECT 3.1950 0.8625 3.3150 1.1250 ;
        RECT 1.8375 0.9750 3.1950 1.1250 ;
        RECT 1.7325 0.7500 1.8375 1.1250 ;
        RECT 1.4025 0.9750 1.7325 1.1250 ;
        RECT 1.2975 0.8325 1.4025 1.1250 ;
        RECT 0.3675 0.9750 1.2975 1.1250 ;
        RECT 0.2625 0.8250 0.3675 1.1250 ;
        RECT 0.0000 0.9750 0.2625 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 4.0650 0.2175 4.1250 0.2775 ;
        RECT 4.0650 0.7800 4.1250 0.8400 ;
        RECT 3.9525 0.4650 4.0125 0.5250 ;
        RECT 3.8550 0.2250 3.9150 0.2850 ;
        RECT 3.8550 0.6525 3.9150 0.7125 ;
        RECT 3.7500 0.4650 3.8100 0.5250 ;
        RECT 3.6450 0.1275 3.7050 0.1875 ;
        RECT 3.6450 0.8325 3.7050 0.8925 ;
        RECT 3.5400 0.4650 3.6000 0.5250 ;
        RECT 3.4350 0.2250 3.4950 0.2850 ;
        RECT 3.4350 0.6525 3.4950 0.7125 ;
        RECT 3.3300 0.4650 3.3900 0.5250 ;
        RECT 3.2250 0.2025 3.2850 0.2625 ;
        RECT 3.2250 0.8700 3.2850 0.9300 ;
        RECT 3.1200 0.4800 3.1800 0.5400 ;
        RECT 3.0150 0.1800 3.0750 0.2400 ;
        RECT 3.0150 0.8100 3.0750 0.8700 ;
        RECT 2.9100 0.4800 2.9700 0.5400 ;
        RECT 2.8050 0.1725 2.8650 0.2325 ;
        RECT 2.8050 0.8250 2.8650 0.8850 ;
        RECT 2.6925 0.4950 2.7525 0.5550 ;
        RECT 2.5950 0.1875 2.6550 0.2475 ;
        RECT 2.5950 0.8175 2.6550 0.8775 ;
        RECT 2.4900 0.6450 2.5500 0.7050 ;
        RECT 2.3850 0.2400 2.4450 0.3000 ;
        RECT 2.3850 0.8175 2.4450 0.8775 ;
        RECT 2.2800 0.4950 2.3400 0.5550 ;
        RECT 2.1750 0.1200 2.2350 0.1800 ;
        RECT 2.0700 0.4950 2.1300 0.5550 ;
        RECT 1.9650 0.2475 2.0250 0.3075 ;
        RECT 1.9650 0.7575 2.0250 0.8175 ;
        RECT 1.8600 0.4800 1.9200 0.5400 ;
        RECT 1.7550 0.7725 1.8150 0.8325 ;
        RECT 1.6500 0.4800 1.7100 0.5400 ;
        RECT 1.5450 0.2550 1.6050 0.3150 ;
        RECT 1.5450 0.8175 1.6050 0.8775 ;
        RECT 1.4475 0.4800 1.5075 0.5400 ;
        RECT 1.3350 0.2250 1.3950 0.2850 ;
        RECT 1.3350 0.8625 1.3950 0.9225 ;
        RECT 1.2300 0.4800 1.2900 0.5400 ;
        RECT 1.1250 0.1800 1.1850 0.2400 ;
        RECT 1.1250 0.7200 1.1850 0.7800 ;
        RECT 1.0200 0.4950 1.0800 0.5550 ;
        RECT 0.9150 0.1725 0.9750 0.2325 ;
        RECT 0.9150 0.8325 0.9750 0.8925 ;
        RECT 0.8100 0.3525 0.8700 0.4125 ;
        RECT 0.7050 0.1650 0.7650 0.2250 ;
        RECT 0.7050 0.8325 0.7650 0.8925 ;
        RECT 0.6000 0.6600 0.6600 0.7200 ;
        RECT 0.3900 0.4200 0.4500 0.4800 ;
        RECT 0.3900 0.6600 0.4500 0.7200 ;
        RECT 0.2850 0.1575 0.3450 0.2175 ;
        RECT 0.2850 0.8475 0.3450 0.9075 ;
        RECT 0.1875 0.5175 0.2475 0.5775 ;
        RECT 0.0750 0.2700 0.1350 0.3300 ;
        RECT 0.0750 0.8175 0.1350 0.8775 ;
        LAYER M1 ;
        RECT 3.9900 0.4425 4.0950 0.6825 ;
        RECT 3.2925 0.4425 3.9900 0.5475 ;
        RECT 3.8325 0.1950 3.9150 0.3675 ;
        RECT 3.4350 0.6225 3.9150 0.7425 ;
        RECT 3.5175 0.2775 3.8325 0.3675 ;
        RECT 3.4125 0.1950 3.5175 0.3675 ;
        RECT 3.2175 0.6450 3.3375 0.7875 ;
        RECT 3.1725 0.4650 3.2175 0.7875 ;
        RECT 3.1425 0.4650 3.1725 0.7050 ;
        RECT 3.0450 0.1500 3.1500 0.3900 ;
        RECT 3.0900 0.4650 3.1425 0.5700 ;
        RECT 3.0675 0.7800 3.0975 0.9000 ;
        RECT 2.9925 0.6450 3.0675 0.9000 ;
        RECT 2.7825 0.1500 3.0450 0.2550 ;
        RECT 2.9700 0.4650 3.0150 0.5700 ;
        RECT 2.4600 0.6450 2.9925 0.7200 ;
        RECT 2.8875 0.3300 2.9700 0.5700 ;
        RECT 2.5425 0.7950 2.9175 0.9000 ;
        RECT 2.7825 0.3300 2.8875 0.4050 ;
        RECT 2.5875 0.4800 2.7825 0.5700 ;
        RECT 2.6550 0.1500 2.6775 0.2850 ;
        RECT 2.5275 0.1500 2.6550 0.3900 ;
        RECT 2.4300 0.4650 2.5875 0.5700 ;
        RECT 2.3475 0.7950 2.4675 0.9000 ;
        RECT 2.3775 0.1950 2.4525 0.3375 ;
        RECT 2.0400 0.2625 2.3775 0.3375 ;
        RECT 2.1300 0.4125 2.3550 0.5850 ;
        RECT 2.2050 0.6600 2.3475 0.9000 ;
        RECT 2.0550 0.4125 2.1300 0.8400 ;
        RECT 1.9425 0.7350 2.0550 0.8400 ;
        RECT 1.9500 0.2175 2.0400 0.3375 ;
        RECT 1.4475 0.4500 1.9500 0.5700 ;
        RECT 1.5150 0.2025 1.8225 0.3750 ;
        RECT 1.4925 0.6600 1.6575 0.9000 ;
        RECT 1.2675 0.4575 1.3725 0.7575 ;
        RECT 1.1925 0.4575 1.2675 0.5925 ;
        RECT 1.0500 0.1500 1.2150 0.3825 ;
        RECT 1.1175 0.6675 1.1925 0.8325 ;
        RECT 0.6900 0.6675 1.1175 0.7425 ;
        RECT 1.0050 0.4875 1.1100 0.5925 ;
        RECT 0.8850 0.1500 1.0500 0.2550 ;
        RECT 0.4575 0.4875 1.0050 0.5625 ;
        RECT 0.5850 0.8175 1.0050 0.9000 ;
        RECT 0.5625 0.3300 0.9450 0.4125 ;
        RECT 0.4650 0.1500 0.7950 0.2550 ;
        RECT 0.5775 0.6375 0.6900 0.7425 ;
        RECT 0.3675 0.6375 0.4800 0.7425 ;
        RECT 0.3825 0.3375 0.4575 0.5625 ;
        RECT 0.1425 0.3375 0.3825 0.4125 ;
        RECT 0.3075 0.6375 0.3675 0.7200 ;
        RECT 0.2325 0.4875 0.3075 0.7200 ;
        RECT 0.1875 0.4875 0.2325 0.6075 ;
        RECT 0.1125 0.7950 0.1575 0.9000 ;
        RECT 0.1125 0.2400 0.1425 0.4125 ;
        RECT 0.0375 0.2400 0.1125 0.9000 ;
        LAYER VIA1 ;
        RECT 3.9900 0.5625 4.0650 0.6375 ;
        RECT 3.3300 0.4575 3.4050 0.5325 ;
        RECT 3.0600 0.2775 3.1350 0.3525 ;
        RECT 2.8275 0.3300 2.9025 0.4050 ;
        RECT 2.7525 0.6450 2.8275 0.7200 ;
        RECT 2.5800 0.8100 2.6550 0.8850 ;
        RECT 2.5650 0.1650 2.6400 0.2400 ;
        RECT 2.4675 0.4800 2.5425 0.5550 ;
        RECT 2.2350 0.7125 2.3100 0.7875 ;
        RECT 2.1225 0.4125 2.1975 0.4875 ;
        RECT 1.8000 0.4650 1.8750 0.5400 ;
        RECT 1.7325 0.2625 1.8075 0.3375 ;
        RECT 1.5375 0.7125 1.6125 0.7875 ;
        RECT 1.1175 0.7125 1.1925 0.7875 ;
        RECT 1.0950 0.2925 1.1700 0.3675 ;
        RECT 0.8550 0.8175 0.9300 0.8925 ;
        RECT 0.5100 0.1650 0.5850 0.2400 ;
        LAYER M2 ;
        RECT 3.9975 0.5625 4.1400 0.6375 ;
        RECT 3.9225 0.5625 3.9975 0.9375 ;
        RECT 2.6550 0.8625 3.9225 0.9375 ;
        RECT 3.3225 0.4200 3.4200 0.5700 ;
        RECT 3.2475 0.1125 3.3225 0.5700 ;
        RECT 2.7000 0.1125 3.2475 0.1875 ;
        RECT 3.0675 0.2625 3.1725 0.3675 ;
        RECT 2.9925 0.2625 3.0675 0.6375 ;
        RECT 2.8425 0.5625 2.9925 0.6375 ;
        RECT 2.8125 0.2925 2.9175 0.4425 ;
        RECT 2.7375 0.5625 2.8425 0.7650 ;
        RECT 2.2725 0.3150 2.8125 0.3900 ;
        RECT 2.6250 0.1125 2.7000 0.2400 ;
        RECT 2.5800 0.7650 2.6550 0.9375 ;
        RECT 2.4900 0.1650 2.6250 0.2400 ;
        RECT 2.4375 0.4650 2.5800 0.5700 ;
        RECT 2.3475 0.4650 2.4375 0.6375 ;
        RECT 1.4625 0.7125 2.3850 0.7875 ;
        RECT 1.8750 0.5625 2.3475 0.6375 ;
        RECT 2.1975 0.3150 2.2725 0.4875 ;
        RECT 2.0250 0.4125 2.1975 0.4875 ;
        RECT 1.9500 0.2625 2.0250 0.4875 ;
        RECT 1.6575 0.2625 1.9500 0.3375 ;
        RECT 1.8000 0.4125 1.8750 0.6375 ;
        RECT 1.5075 0.4125 1.8000 0.4875 ;
        RECT 1.4325 0.1350 1.5075 0.4875 ;
        RECT 0.9450 0.1350 1.4325 0.2100 ;
        RECT 1.0950 0.7125 1.2675 0.7875 ;
        RECT 1.0950 0.2925 1.2450 0.3675 ;
        RECT 1.0200 0.2925 1.0950 0.7875 ;
        RECT 0.8700 0.1350 0.9450 0.9300 ;
        RECT 0.4350 0.1650 0.8700 0.2400 ;
        RECT 0.8400 0.7800 0.8700 0.9300 ;
    END
END XNR3_0111


MACRO XNR3_1000
    CLASS CORE ;
    FOREIGN XNR3_1000 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.7700 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 7.0875 0.3075 7.4025 0.7425 ;
        VIA 7.2450 0.3750 VIA12_slot ;
        VIA 7.2450 0.6750 VIA12_slot ;
        END
    END ZN
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 5.5425 0.4125 6.0975 0.4875 ;
        RECT 5.4375 0.4125 5.5425 0.6075 ;
        VIA 5.9775 0.4500 VIA12_square ;
        VIA 5.4900 0.5175 VIA12_square ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.9000 0.4350 1.0125 0.6375 ;
        RECT 0.3900 0.5625 0.9000 0.6375 ;
        VIA 0.9600 0.5175 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 2.1825 0.4125 2.7375 0.4875 ;
        RECT 2.0775 0.4125 2.1825 0.6075 ;
        VIA 2.6175 0.4500 VIA12_square ;
        VIA 2.1300 0.5175 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 5.8500 -0.0750 7.7700 0.0750 ;
        RECT 5.7000 -0.0750 5.8500 0.2175 ;
        RECT 5.4150 -0.0750 5.7000 0.0750 ;
        RECT 5.2950 -0.0750 5.4150 0.2250 ;
        RECT 4.9950 -0.0750 5.2950 0.0750 ;
        RECT 4.8750 -0.0750 4.9950 0.2325 ;
        RECT 4.5750 -0.0750 4.8750 0.0750 ;
        RECT 4.4550 -0.0750 4.5750 0.2325 ;
        RECT 2.4900 -0.0750 4.4550 0.0750 ;
        RECT 2.3400 -0.0750 2.4900 0.2175 ;
        RECT 2.0550 -0.0750 2.3400 0.0750 ;
        RECT 1.9350 -0.0750 2.0550 0.2250 ;
        RECT 1.6350 -0.0750 1.9350 0.0750 ;
        RECT 1.5150 -0.0750 1.6350 0.2325 ;
        RECT 1.2150 -0.0750 1.5150 0.0750 ;
        RECT 1.0950 -0.0750 1.2150 0.2325 ;
        RECT 0.7950 -0.0750 1.0950 0.0750 ;
        RECT 0.6750 -0.0750 0.7950 0.2325 ;
        RECT 0.3675 -0.0750 0.6750 0.0750 ;
        RECT 0.2625 -0.0750 0.3675 0.2325 ;
        RECT 0.0000 -0.0750 0.2625 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 5.8350 0.9750 7.7700 1.1250 ;
        RECT 5.7150 0.8325 5.8350 1.1250 ;
        RECT 5.4300 0.9750 5.7150 1.1250 ;
        RECT 5.2800 0.8325 5.4300 1.1250 ;
        RECT 4.9950 0.9750 5.2800 1.1250 ;
        RECT 4.8750 0.8400 4.9950 1.1250 ;
        RECT 4.5750 0.9750 4.8750 1.1250 ;
        RECT 4.4550 0.8250 4.5750 1.1250 ;
        RECT 2.4750 0.9750 4.4550 1.1250 ;
        RECT 2.3550 0.8325 2.4750 1.1250 ;
        RECT 2.0700 0.9750 2.3550 1.1250 ;
        RECT 1.9200 0.8325 2.0700 1.1250 ;
        RECT 1.6350 0.9750 1.9200 1.1250 ;
        RECT 1.5150 0.8400 1.6350 1.1250 ;
        RECT 1.2150 0.9750 1.5150 1.1250 ;
        RECT 1.0950 0.8400 1.2150 1.1250 ;
        RECT 0.7950 0.9750 1.0950 1.1250 ;
        RECT 0.6750 0.8400 0.7950 1.1250 ;
        RECT 0.3750 0.9750 0.6750 1.1250 ;
        RECT 0.2550 0.8400 0.3750 1.1250 ;
        RECT 0.0000 0.9750 0.2550 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 7.6350 0.3075 7.6950 0.3675 ;
        RECT 7.6350 0.6750 7.6950 0.7350 ;
        RECT 7.5300 0.4950 7.5900 0.5550 ;
        RECT 7.4250 0.1575 7.4850 0.2175 ;
        RECT 7.4250 0.8325 7.4850 0.8925 ;
        RECT 7.3200 0.4950 7.3800 0.5550 ;
        RECT 7.2150 0.3225 7.2750 0.3825 ;
        RECT 7.2150 0.6750 7.2750 0.7350 ;
        RECT 7.1100 0.4950 7.1700 0.5550 ;
        RECT 7.0050 0.1575 7.0650 0.2175 ;
        RECT 7.0050 0.8325 7.0650 0.8925 ;
        RECT 6.9000 0.4950 6.9600 0.5550 ;
        RECT 6.7950 0.2625 6.8550 0.3225 ;
        RECT 6.7950 0.6750 6.8550 0.7350 ;
        RECT 6.6900 0.4800 6.7500 0.5400 ;
        RECT 6.5850 0.3000 6.6450 0.3600 ;
        RECT 6.5850 0.6675 6.6450 0.7275 ;
        RECT 6.4800 0.4800 6.5400 0.5400 ;
        RECT 6.3750 0.1575 6.4350 0.2175 ;
        RECT 6.3750 0.8325 6.4350 0.8925 ;
        RECT 6.2700 0.4800 6.3300 0.5400 ;
        RECT 6.1650 0.3000 6.2250 0.3600 ;
        RECT 6.1650 0.6825 6.2250 0.7425 ;
        RECT 6.0600 0.4800 6.1200 0.5400 ;
        RECT 5.9550 0.1875 6.0150 0.2475 ;
        RECT 5.9550 0.8025 6.0150 0.8625 ;
        RECT 5.7450 0.1575 5.8050 0.2175 ;
        RECT 5.7450 0.8325 5.8050 0.8925 ;
        RECT 5.6400 0.4875 5.7000 0.5475 ;
        RECT 5.5350 0.3075 5.5950 0.3675 ;
        RECT 5.5350 0.6900 5.5950 0.7500 ;
        RECT 5.4300 0.4875 5.4900 0.5475 ;
        RECT 5.3250 0.1425 5.3850 0.2025 ;
        RECT 5.3250 0.8325 5.3850 0.8925 ;
        RECT 5.2200 0.4875 5.2800 0.5475 ;
        RECT 5.1150 0.2925 5.1750 0.3525 ;
        RECT 5.1150 0.7200 5.1750 0.7800 ;
        RECT 5.0100 0.4875 5.0700 0.5475 ;
        RECT 4.9050 0.1650 4.9650 0.2250 ;
        RECT 4.9050 0.8475 4.9650 0.9075 ;
        RECT 4.8000 0.4875 4.8600 0.5475 ;
        RECT 4.6950 0.2925 4.7550 0.3525 ;
        RECT 4.6950 0.7350 4.7550 0.7950 ;
        RECT 4.5900 0.4875 4.6500 0.5475 ;
        RECT 4.4850 0.1650 4.5450 0.2250 ;
        RECT 4.4850 0.8325 4.5450 0.8925 ;
        RECT 4.2750 0.3075 4.3350 0.3675 ;
        RECT 4.2750 0.6750 4.3350 0.7350 ;
        RECT 4.1700 0.4950 4.2300 0.5550 ;
        RECT 4.0650 0.1575 4.1250 0.2175 ;
        RECT 4.0650 0.8325 4.1250 0.8925 ;
        RECT 3.9600 0.4950 4.0200 0.5550 ;
        RECT 3.8550 0.3225 3.9150 0.3825 ;
        RECT 3.8550 0.6750 3.9150 0.7350 ;
        RECT 3.7500 0.4950 3.8100 0.5550 ;
        RECT 3.6450 0.1575 3.7050 0.2175 ;
        RECT 3.6450 0.8325 3.7050 0.8925 ;
        RECT 3.5400 0.4950 3.6000 0.5550 ;
        RECT 3.4350 0.2625 3.4950 0.3225 ;
        RECT 3.4350 0.6750 3.4950 0.7350 ;
        RECT 3.3300 0.4800 3.3900 0.5400 ;
        RECT 3.2250 0.3000 3.2850 0.3600 ;
        RECT 3.2250 0.6675 3.2850 0.7275 ;
        RECT 3.1200 0.4800 3.1800 0.5400 ;
        RECT 3.0150 0.1575 3.0750 0.2175 ;
        RECT 3.0150 0.8325 3.0750 0.8925 ;
        RECT 2.9100 0.4800 2.9700 0.5400 ;
        RECT 2.8050 0.3000 2.8650 0.3600 ;
        RECT 2.8050 0.6825 2.8650 0.7425 ;
        RECT 2.7000 0.4800 2.7600 0.5400 ;
        RECT 2.5950 0.1875 2.6550 0.2475 ;
        RECT 2.5950 0.8025 2.6550 0.8625 ;
        RECT 2.3850 0.1575 2.4450 0.2175 ;
        RECT 2.3850 0.8325 2.4450 0.8925 ;
        RECT 2.2800 0.4875 2.3400 0.5475 ;
        RECT 2.1750 0.3075 2.2350 0.3675 ;
        RECT 2.1750 0.6900 2.2350 0.7500 ;
        RECT 2.0700 0.4875 2.1300 0.5475 ;
        RECT 1.9650 0.1425 2.0250 0.2025 ;
        RECT 1.9650 0.8325 2.0250 0.8925 ;
        RECT 1.8600 0.4875 1.9200 0.5475 ;
        RECT 1.7550 0.2925 1.8150 0.3525 ;
        RECT 1.7550 0.7200 1.8150 0.7800 ;
        RECT 1.6500 0.4875 1.7100 0.5475 ;
        RECT 1.5450 0.1650 1.6050 0.2250 ;
        RECT 1.5450 0.8475 1.6050 0.9075 ;
        RECT 1.4400 0.4875 1.5000 0.5475 ;
        RECT 1.3350 0.2925 1.3950 0.3525 ;
        RECT 1.3350 0.7350 1.3950 0.7950 ;
        RECT 1.2300 0.4875 1.2900 0.5475 ;
        RECT 1.1250 0.1650 1.1850 0.2250 ;
        RECT 1.1250 0.8475 1.1850 0.9075 ;
        RECT 1.0200 0.4875 1.0800 0.5475 ;
        RECT 0.9150 0.2925 0.9750 0.3525 ;
        RECT 0.9150 0.7350 0.9750 0.7950 ;
        RECT 0.8100 0.4875 0.8700 0.5475 ;
        RECT 0.7050 0.1650 0.7650 0.2250 ;
        RECT 0.7050 0.8475 0.7650 0.9075 ;
        RECT 0.6000 0.4875 0.6600 0.5475 ;
        RECT 0.4950 0.2925 0.5550 0.3525 ;
        RECT 0.4950 0.7350 0.5550 0.7950 ;
        RECT 0.3900 0.4875 0.4500 0.5475 ;
        RECT 0.2850 0.1500 0.3450 0.2100 ;
        RECT 0.2850 0.8475 0.3450 0.9075 ;
        RECT 0.1800 0.4875 0.2400 0.5475 ;
        RECT 0.0750 0.2925 0.1350 0.3525 ;
        RECT 0.0750 0.7350 0.1350 0.7950 ;
        LAYER M1 ;
        RECT 7.6050 0.2775 7.7250 0.4125 ;
        RECT 7.6200 0.6375 7.7025 0.7875 ;
        RECT 7.0200 0.4875 7.6500 0.5625 ;
        RECT 7.0875 0.6375 7.6200 0.7350 ;
        RECT 7.0875 0.3075 7.6050 0.4125 ;
        RECT 7.1325 0.1500 7.5375 0.2250 ;
        RECT 7.0875 0.8250 7.5150 0.9000 ;
        RECT 6.9675 0.1500 7.1325 0.2325 ;
        RECT 6.8625 0.3075 7.0875 0.3825 ;
        RECT 6.8175 0.6600 7.0875 0.7350 ;
        RECT 6.9225 0.8175 7.0875 0.9000 ;
        RECT 6.8250 0.4575 7.0200 0.5850 ;
        RECT 6.7875 0.1500 6.8625 0.3825 ;
        RECT 6.7425 0.6600 6.8175 0.9000 ;
        RECT 6.0300 0.1500 6.7875 0.2250 ;
        RECT 6.6450 0.4500 6.7500 0.5700 ;
        RECT 6.0225 0.8250 6.7425 0.9000 ;
        RECT 6.1350 0.3000 6.6750 0.3750 ;
        RECT 6.5025 0.6450 6.6675 0.7500 ;
        RECT 6.0300 0.4500 6.6450 0.5400 ;
        RECT 6.1350 0.6750 6.5025 0.7500 ;
        RECT 5.9250 0.1500 6.0300 0.2850 ;
        RECT 5.9250 0.3750 6.0300 0.5400 ;
        RECT 5.9475 0.7575 6.0225 0.9000 ;
        RECT 5.7750 0.3075 5.8500 0.7575 ;
        RECT 5.4975 0.3075 5.7750 0.3825 ;
        RECT 5.4300 0.6525 5.7750 0.7575 ;
        RECT 5.3925 0.4575 5.7000 0.5775 ;
        RECT 5.1825 0.3075 5.3100 0.3825 ;
        RECT 4.5300 0.4725 5.3100 0.5775 ;
        RECT 5.0925 0.2625 5.1825 0.3825 ;
        RECT 5.1075 0.6675 5.1825 0.8175 ;
        RECT 4.7625 0.6675 5.1075 0.7425 ;
        RECT 4.7775 0.3075 5.0925 0.3825 ;
        RECT 4.6725 0.2625 4.7775 0.3825 ;
        RECT 4.6875 0.6675 4.7625 0.8400 ;
        RECT 4.4550 0.3075 4.5300 0.7350 ;
        RECT 3.5025 0.3075 4.4550 0.3825 ;
        RECT 3.4575 0.6600 4.4550 0.7350 ;
        RECT 3.6600 0.4875 4.2900 0.5625 ;
        RECT 3.7725 0.1500 4.1775 0.2250 ;
        RECT 3.7275 0.8250 4.1550 0.9000 ;
        RECT 3.6075 0.1500 3.7725 0.2325 ;
        RECT 3.5625 0.8175 3.7275 0.9000 ;
        RECT 3.4650 0.4575 3.6600 0.5850 ;
        RECT 3.4275 0.1500 3.5025 0.3825 ;
        RECT 3.3825 0.6600 3.4575 0.9000 ;
        RECT 2.6700 0.1500 3.4275 0.2250 ;
        RECT 3.2850 0.4500 3.3900 0.5700 ;
        RECT 2.6625 0.8250 3.3825 0.9000 ;
        RECT 2.7750 0.3000 3.3150 0.3750 ;
        RECT 3.1425 0.6450 3.3075 0.7500 ;
        RECT 2.6700 0.4500 3.2850 0.5400 ;
        RECT 2.7750 0.6750 3.1425 0.7500 ;
        RECT 2.5650 0.1500 2.6700 0.2850 ;
        RECT 2.5650 0.3750 2.6700 0.5400 ;
        RECT 2.5875 0.7575 2.6625 0.9000 ;
        RECT 2.4150 0.3075 2.4900 0.7575 ;
        RECT 2.1375 0.3075 2.4150 0.3825 ;
        RECT 2.0700 0.6525 2.4150 0.7575 ;
        RECT 2.0325 0.4575 2.3400 0.5775 ;
        RECT 1.8225 0.3000 2.0250 0.3825 ;
        RECT 1.7925 0.4725 1.9500 0.5775 ;
        RECT 1.7475 0.2625 1.8225 0.3825 ;
        RECT 1.7475 0.6825 1.8225 0.8175 ;
        RECT 1.2300 0.4575 1.7925 0.5775 ;
        RECT 1.4025 0.3075 1.7475 0.3825 ;
        RECT 1.4025 0.6825 1.7475 0.7575 ;
        RECT 1.3275 0.2250 1.4025 0.3825 ;
        RECT 1.3275 0.6825 1.4025 0.8400 ;
        RECT 1.1550 0.3075 1.2300 0.7575 ;
        RECT 0.9825 0.3075 1.1550 0.3825 ;
        RECT 0.9825 0.6825 1.1550 0.7575 ;
        RECT 0.1500 0.4575 1.0800 0.5775 ;
        RECT 0.9075 0.2325 0.9825 0.3825 ;
        RECT 0.9075 0.6825 0.9825 0.8400 ;
        RECT 0.5625 0.3075 0.9075 0.3825 ;
        RECT 0.5625 0.6825 0.9075 0.7575 ;
        RECT 0.4875 0.2325 0.5625 0.3825 ;
        RECT 0.4875 0.6825 0.5625 0.8400 ;
        RECT 0.1425 0.3075 0.4875 0.3825 ;
        RECT 0.1425 0.6825 0.4875 0.7575 ;
        RECT 0.0675 0.2325 0.1425 0.3825 ;
        RECT 0.0675 0.6825 0.1425 0.8400 ;
        LAYER VIA1 ;
        RECT 7.0125 0.1575 7.0875 0.2325 ;
        RECT 6.9675 0.8175 7.0425 0.8925 ;
        RECT 6.8625 0.4800 6.9375 0.5550 ;
        RECT 6.5475 0.6675 6.6225 0.7425 ;
        RECT 6.3225 0.3000 6.3975 0.3750 ;
        RECT 5.7750 0.5625 5.8500 0.6375 ;
        RECT 5.1675 0.3075 5.2425 0.3825 ;
        RECT 4.9800 0.4875 5.0550 0.5625 ;
        RECT 4.8300 0.6675 4.9050 0.7425 ;
        RECT 4.7850 0.3075 4.8600 0.3825 ;
        RECT 3.6525 0.1575 3.7275 0.2325 ;
        RECT 3.6075 0.8175 3.6825 0.8925 ;
        RECT 3.5175 0.4800 3.5925 0.5550 ;
        RECT 3.1875 0.6675 3.2625 0.7425 ;
        RECT 2.9625 0.3000 3.0375 0.3750 ;
        RECT 2.4150 0.5625 2.4900 0.6375 ;
        RECT 1.9050 0.3075 1.9800 0.3825 ;
        RECT 1.7475 0.4875 1.8225 0.5625 ;
        RECT 1.5375 0.6825 1.6125 0.7575 ;
        RECT 1.4625 0.3075 1.5375 0.3825 ;
        LAYER M2 ;
        RECT 6.9675 0.1125 7.1325 0.2325 ;
        RECT 6.9225 0.8175 7.0875 0.9375 ;
        RECT 5.0550 0.1125 6.9675 0.1875 ;
        RECT 6.8625 0.4275 6.9375 0.6225 ;
        RECT 4.9050 0.8625 6.9225 0.9375 ;
        RECT 6.6375 0.4275 6.8625 0.5025 ;
        RECT 6.5325 0.6225 6.6450 0.7875 ;
        RECT 6.5625 0.4275 6.6375 0.5475 ;
        RECT 6.4575 0.4725 6.5625 0.5475 ;
        RECT 5.0550 0.7125 6.5325 0.7875 ;
        RECT 6.3825 0.4725 6.4575 0.6375 ;
        RECT 6.2775 0.2625 6.4425 0.3900 ;
        RECT 5.7150 0.5625 6.3825 0.6375 ;
        RECT 5.2575 0.2625 6.2775 0.3375 ;
        RECT 5.1525 0.2625 5.2575 0.4425 ;
        RECT 4.9800 0.1125 5.0550 0.7875 ;
        RECT 4.8300 0.3075 4.9050 0.9375 ;
        RECT 4.7400 0.3075 4.8300 0.3825 ;
        RECT 3.7425 0.1575 3.8250 0.7200 ;
        RECT 3.6075 0.1575 3.7425 0.2325 ;
        RECT 3.3000 0.6450 3.7425 0.7200 ;
        RECT 3.5550 0.8175 3.7275 0.8925 ;
        RECT 3.4650 0.4275 3.6525 0.5700 ;
        RECT 3.4800 0.8175 3.5550 0.9375 ;
        RECT 1.6125 0.8625 3.4800 0.9375 ;
        RECT 3.2775 0.4275 3.4650 0.5025 ;
        RECT 3.1725 0.6225 3.3000 0.7875 ;
        RECT 3.2025 0.4275 3.2775 0.5475 ;
        RECT 3.0975 0.4725 3.2025 0.5475 ;
        RECT 1.8225 0.7125 3.1725 0.7875 ;
        RECT 3.0225 0.4725 3.0975 0.6375 ;
        RECT 2.9175 0.2625 3.0825 0.3900 ;
        RECT 2.3550 0.5625 3.0225 0.6375 ;
        RECT 1.9800 0.2625 2.9175 0.3375 ;
        RECT 1.9050 0.2625 1.9800 0.4500 ;
        RECT 1.7475 0.4125 1.8225 0.7875 ;
        RECT 1.5375 0.3075 1.6125 0.9375 ;
        RECT 1.3875 0.3075 1.5375 0.3825 ;
    END
END XNR3_1000


MACRO XNR3_1010
    CLASS CORE ;
    FOREIGN XNR3_1010 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.1500 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 3.0375 0.1500 3.1125 0.9000 ;
        RECT 2.9850 0.1500 3.0375 0.3825 ;
        RECT 2.9925 0.6675 3.0375 0.9000 ;
        END
    END ZN
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 2.7750 0.1125 3.0900 0.1875 ;
        RECT 2.7000 0.1125 2.7750 0.4875 ;
        RECT 2.3850 0.4125 2.7000 0.4875 ;
        VIA 2.6850 0.4500 VIA12_square ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.2150 0.5625 1.6800 0.6375 ;
        VIA 1.3575 0.6000 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.6075 0.3375 0.7800 0.4425 ;
        RECT 0.5325 0.3375 0.6075 0.6375 ;
        RECT 0.0675 0.5625 0.5325 0.6375 ;
        VIA 0.6975 0.3750 VIA12_square ;
        VIA 0.2700 0.6000 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 2.8950 -0.0750 3.1500 0.0750 ;
        RECT 2.7750 -0.0750 2.8950 0.2550 ;
        RECT 1.8450 -0.0750 2.7750 0.0750 ;
        RECT 1.7250 -0.0750 1.8450 0.2400 ;
        RECT 1.4100 -0.0750 1.7250 0.0750 ;
        RECT 1.3200 -0.0750 1.4100 0.2475 ;
        RECT 0.3675 -0.0750 1.3200 0.0750 ;
        RECT 0.2625 -0.0750 0.3675 0.2475 ;
        RECT 0.0000 -0.0750 0.2625 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 2.8950 0.9750 3.1500 1.1250 ;
        RECT 2.7750 0.8625 2.8950 1.1250 ;
        RECT 1.8450 0.9750 2.7750 1.1250 ;
        RECT 1.7250 0.8250 1.8450 1.1250 ;
        RECT 1.4025 0.9750 1.7250 1.1250 ;
        RECT 1.3275 0.7875 1.4025 1.1250 ;
        RECT 0.3675 0.9750 1.3275 1.1250 ;
        RECT 0.2625 0.8250 0.3675 1.1250 ;
        RECT 0.0000 0.9750 0.2625 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 3.0150 0.1575 3.0750 0.2175 ;
        RECT 3.0150 0.8175 3.0750 0.8775 ;
        RECT 2.9025 0.4875 2.9625 0.5475 ;
        RECT 2.8050 0.1650 2.8650 0.2250 ;
        RECT 2.8050 0.8700 2.8650 0.9300 ;
        RECT 2.7000 0.4650 2.7600 0.5250 ;
        RECT 2.5950 0.1575 2.6550 0.2175 ;
        RECT 2.5950 0.7950 2.6550 0.8550 ;
        RECT 2.4900 0.4500 2.5500 0.5100 ;
        RECT 2.3850 0.1575 2.4450 0.2175 ;
        RECT 2.3850 0.8325 2.4450 0.8925 ;
        RECT 2.2800 0.5025 2.3400 0.5625 ;
        RECT 2.1750 0.1800 2.2350 0.2400 ;
        RECT 2.1750 0.8325 2.2350 0.8925 ;
        RECT 2.0700 0.6600 2.1300 0.7200 ;
        RECT 1.8600 0.3600 1.9200 0.4200 ;
        RECT 1.8600 0.6300 1.9200 0.6900 ;
        RECT 1.7550 0.1575 1.8150 0.2175 ;
        RECT 1.7550 0.8550 1.8150 0.9150 ;
        RECT 1.6500 0.5250 1.7100 0.5850 ;
        RECT 1.5450 0.1575 1.6050 0.2175 ;
        RECT 1.5450 0.8175 1.6050 0.8775 ;
        RECT 1.3350 0.1575 1.3950 0.2175 ;
        RECT 1.3350 0.8175 1.3950 0.8775 ;
        RECT 1.2300 0.5100 1.2900 0.5700 ;
        RECT 1.1250 0.2250 1.1850 0.2850 ;
        RECT 1.1250 0.7350 1.1850 0.7950 ;
        RECT 1.0200 0.4950 1.0800 0.5550 ;
        RECT 0.9150 0.1575 0.9750 0.2175 ;
        RECT 0.9150 0.8325 0.9750 0.8925 ;
        RECT 0.8100 0.3525 0.8700 0.4125 ;
        RECT 0.7050 0.1650 0.7650 0.2250 ;
        RECT 0.7050 0.8325 0.7650 0.8925 ;
        RECT 0.6000 0.6600 0.6600 0.7200 ;
        RECT 0.3900 0.4200 0.4500 0.4800 ;
        RECT 0.3900 0.6600 0.4500 0.7200 ;
        RECT 0.2850 0.1575 0.3450 0.2175 ;
        RECT 0.2850 0.8475 0.3450 0.9075 ;
        RECT 0.1875 0.5175 0.2475 0.5775 ;
        RECT 0.0750 0.1575 0.1350 0.2175 ;
        RECT 0.0750 0.8175 0.1350 0.8775 ;
        LAYER M1 ;
        RECT 2.9175 0.4575 2.9625 0.5775 ;
        RECT 2.8425 0.4575 2.9175 0.7875 ;
        RECT 2.7675 0.6825 2.8425 0.7875 ;
        RECT 2.6325 0.3300 2.7675 0.5700 ;
        RECT 2.4825 0.1500 2.6925 0.2550 ;
        RECT 2.5800 0.6450 2.6850 0.8850 ;
        RECT 2.0400 0.6450 2.5800 0.7350 ;
        RECT 2.4825 0.3450 2.5575 0.5400 ;
        RECT 2.3100 0.1500 2.4825 0.2700 ;
        RECT 1.6350 0.3450 2.4825 0.4200 ;
        RECT 2.1000 0.8100 2.4750 0.9000 ;
        RECT 1.9350 0.4950 2.3775 0.5700 ;
        RECT 1.9275 0.1500 2.2350 0.2700 ;
        RECT 1.8300 0.4950 1.9350 0.7200 ;
        RECT 1.6425 0.4950 1.8300 0.6150 ;
        RECT 1.5675 0.1500 1.6350 0.4200 ;
        RECT 1.5675 0.7950 1.6275 0.9000 ;
        RECT 1.5150 0.1500 1.5675 0.9000 ;
        RECT 1.4850 0.3450 1.5150 0.9000 ;
        RECT 1.3050 0.4875 1.4100 0.6825 ;
        RECT 1.1925 0.4875 1.3050 0.5925 ;
        RECT 1.0575 0.1500 1.2150 0.4125 ;
        RECT 1.1100 0.6675 1.2150 0.8325 ;
        RECT 1.0050 0.4875 1.1100 0.5925 ;
        RECT 0.6900 0.6675 1.1100 0.7425 ;
        RECT 0.8850 0.1500 1.0575 0.2550 ;
        RECT 0.4575 0.4875 1.0050 0.5625 ;
        RECT 0.5850 0.8175 1.0050 0.9000 ;
        RECT 0.5625 0.3300 0.9450 0.4125 ;
        RECT 0.4650 0.1500 0.7950 0.2550 ;
        RECT 0.5775 0.6375 0.6900 0.7425 ;
        RECT 0.3675 0.6375 0.4800 0.7425 ;
        RECT 0.3825 0.3375 0.4575 0.5625 ;
        RECT 0.1650 0.3375 0.3825 0.4125 ;
        RECT 0.3075 0.6375 0.3675 0.7200 ;
        RECT 0.2325 0.4875 0.3075 0.7200 ;
        RECT 0.1875 0.4875 0.2325 0.6075 ;
        RECT 0.1125 0.1500 0.1650 0.4125 ;
        RECT 0.1125 0.7950 0.1575 0.9000 ;
        RECT 0.0375 0.1500 0.1125 0.9000 ;
        LAYER VIA1 ;
        RECT 2.8425 0.5625 2.9175 0.6375 ;
        RECT 2.4075 0.6450 2.4825 0.7200 ;
        RECT 2.3475 0.1725 2.4225 0.2475 ;
        RECT 2.2575 0.8100 2.3325 0.8850 ;
        RECT 1.9875 0.1800 2.0625 0.2550 ;
        RECT 1.8375 0.4950 1.9125 0.5700 ;
        RECT 1.0950 0.3225 1.1700 0.3975 ;
        RECT 1.0200 0.6675 1.0950 0.7425 ;
        RECT 0.8250 0.8175 0.9000 0.8925 ;
        RECT 0.5100 0.1725 0.5850 0.2475 ;
        LAYER M2 ;
        RECT 2.7525 0.5625 3.0000 0.6375 ;
        RECT 2.6775 0.5625 2.7525 0.8850 ;
        RECT 2.1150 0.8100 2.6775 0.8850 ;
        RECT 2.2650 0.6450 2.5275 0.7200 ;
        RECT 2.2650 0.1725 2.4675 0.2475 ;
        RECT 2.1900 0.1725 2.2650 0.7200 ;
        RECT 2.0400 0.1650 2.1150 0.8850 ;
        RECT 1.9500 0.1650 2.0400 0.2700 ;
        RECT 1.8375 0.4125 1.9125 0.6450 ;
        RECT 1.4325 0.4125 1.8375 0.4875 ;
        RECT 1.3575 0.1575 1.4325 0.4875 ;
        RECT 0.9450 0.1575 1.3575 0.2325 ;
        RECT 1.0950 0.3075 1.2150 0.4125 ;
        RECT 1.0200 0.3075 1.0950 0.7950 ;
        RECT 0.8700 0.1575 0.9450 0.9000 ;
        RECT 0.6225 0.1575 0.8700 0.2325 ;
        RECT 0.7800 0.8100 0.8700 0.9000 ;
        RECT 0.4725 0.1575 0.6225 0.2625 ;
    END
END XNR3_1010


MACRO XNR4_0111
    CLASS CORE ;
    FOREIGN XNR4_0111 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.3000 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 3.3075 0.2625 3.6225 0.7125 ;
        VIA 3.4650 0.3225 VIA12_slot ;
        VIA 3.4650 0.6525 VIA12_slot ;
        END
    END ZN
    PIN A4
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.5175 0.5625 0.7125 0.6375 ;
        RECT 0.3525 0.4950 0.5175 0.6375 ;
        RECT 0.0675 0.5625 0.3525 0.6375 ;
        VIA 0.4350 0.5400 VIA12_square ;
        END
    END A4
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.3500 0.8625 1.6125 0.9375 ;
        RECT 1.2750 0.5925 1.3500 0.9375 ;
        RECT 1.0725 0.8625 1.2750 0.9375 ;
        VIA 1.3125 0.6750 VIA12_square ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 4.1475 0.4125 4.2825 0.4875 ;
        RECT 4.0425 0.4125 4.1475 0.6075 ;
        RECT 3.7425 0.4125 4.0425 0.4875 ;
        VIA 4.0950 0.5250 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 5.2725 0.4125 6.1575 0.4875 ;
        RECT 5.1975 0.3225 5.2725 0.4875 ;
        RECT 4.7025 0.3225 5.1975 0.4050 ;
        RECT 4.6275 0.3225 4.7025 0.4950 ;
        VIA 6.0450 0.4500 VIA12_square ;
        VIA 5.3625 0.4500 VIA12_square ;
        VIA 4.6650 0.4125 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 6.2475 -0.0750 6.3000 0.0750 ;
        RECT 6.1425 -0.0750 6.2475 0.2850 ;
        RECT 5.4150 -0.0750 6.1425 0.0750 ;
        RECT 5.2950 -0.0750 5.4150 0.1875 ;
        RECT 4.3425 -0.0750 5.2950 0.0750 ;
        RECT 4.2375 -0.0750 4.3425 0.2475 ;
        RECT 3.9225 -0.0750 4.2375 0.0750 ;
        RECT 3.8475 -0.0750 3.9225 0.3150 ;
        RECT 3.5250 -0.0750 3.8475 0.0750 ;
        RECT 3.4050 -0.0750 3.5250 0.2025 ;
        RECT 3.0900 -0.0750 3.4050 0.0750 ;
        RECT 3.0150 -0.0750 3.0900 0.2625 ;
        RECT 2.6550 -0.0750 3.0150 0.0750 ;
        RECT 2.5800 -0.0750 2.6550 0.2625 ;
        RECT 1.4250 -0.0750 2.5800 0.0750 ;
        RECT 1.3050 -0.0750 1.4250 0.2400 ;
        RECT 0.3750 -0.0750 1.3050 0.0750 ;
        RECT 0.2550 -0.0750 0.3750 0.1875 ;
        RECT 0.0000 -0.0750 0.2550 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 6.0450 0.9750 6.3000 1.1250 ;
        RECT 5.9400 0.8100 6.0450 1.1250 ;
        RECT 5.6175 0.9750 5.9400 1.1250 ;
        RECT 5.5125 0.7875 5.6175 1.1250 ;
        RECT 4.3650 0.9750 5.5125 1.1250 ;
        RECT 4.2450 0.8025 4.3650 1.1250 ;
        RECT 3.9450 0.9750 4.2450 1.1250 ;
        RECT 3.8250 0.6525 3.9450 1.1250 ;
        RECT 3.5100 0.9750 3.8250 1.1250 ;
        RECT 3.4200 0.8025 3.5100 1.1250 ;
        RECT 3.0900 0.9750 3.4200 1.1250 ;
        RECT 3.0000 0.7650 3.0900 1.1250 ;
        RECT 2.6850 0.9750 3.0000 1.1250 ;
        RECT 2.5650 0.8700 2.6850 1.1250 ;
        RECT 1.4250 0.9750 2.5650 1.1250 ;
        RECT 1.3050 0.8625 1.4250 1.1250 ;
        RECT 0.3750 0.9750 1.3050 1.1250 ;
        RECT 0.2550 0.8625 0.3750 1.1250 ;
        RECT 0.0000 0.9750 0.2550 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 6.1650 0.2025 6.2250 0.2625 ;
        RECT 6.1650 0.6900 6.2250 0.7500 ;
        RECT 6.0600 0.4725 6.1200 0.5325 ;
        RECT 5.9550 0.1875 6.0150 0.2475 ;
        RECT 5.9550 0.8400 6.0150 0.9000 ;
        RECT 5.8500 0.4800 5.9100 0.5400 ;
        RECT 5.7450 0.8175 5.8050 0.8775 ;
        RECT 5.6400 0.4800 5.7000 0.5400 ;
        RECT 5.5350 0.2700 5.5950 0.3300 ;
        RECT 5.5350 0.8175 5.5950 0.8775 ;
        RECT 5.4300 0.4650 5.4900 0.5250 ;
        RECT 5.3250 0.1275 5.3850 0.1875 ;
        RECT 5.2200 0.4650 5.2800 0.5250 ;
        RECT 5.1150 0.2400 5.1750 0.3000 ;
        RECT 5.1150 0.8175 5.1750 0.8775 ;
        RECT 5.0100 0.6450 5.0700 0.7050 ;
        RECT 4.9050 0.2325 4.9650 0.2925 ;
        RECT 4.9050 0.8175 4.9650 0.8775 ;
        RECT 4.8000 0.4875 4.8600 0.5475 ;
        RECT 4.6950 0.1725 4.7550 0.2325 ;
        RECT 4.6950 0.8250 4.7550 0.8850 ;
        RECT 4.5900 0.4500 4.6500 0.5100 ;
        RECT 4.4850 0.6525 4.5450 0.7125 ;
        RECT 4.2750 0.1575 4.3350 0.2175 ;
        RECT 4.2750 0.8100 4.3350 0.8700 ;
        RECT 4.1700 0.4875 4.2300 0.5475 ;
        RECT 4.0650 0.3075 4.1250 0.3675 ;
        RECT 4.0650 0.7275 4.1250 0.7875 ;
        RECT 3.9600 0.4875 4.0200 0.5475 ;
        RECT 3.8550 0.2250 3.9150 0.2850 ;
        RECT 3.8550 0.6675 3.9150 0.7275 ;
        RECT 3.8550 0.8325 3.9150 0.8925 ;
        RECT 3.7500 0.4650 3.8100 0.5250 ;
        RECT 3.6450 0.2250 3.7050 0.2850 ;
        RECT 3.6450 0.7575 3.7050 0.8175 ;
        RECT 3.5400 0.4650 3.6000 0.5250 ;
        RECT 3.4350 0.1350 3.4950 0.1950 ;
        RECT 3.4350 0.8325 3.4950 0.8925 ;
        RECT 3.3300 0.4650 3.3900 0.5250 ;
        RECT 3.2250 0.2250 3.2850 0.2850 ;
        RECT 3.2250 0.7575 3.2850 0.8175 ;
        RECT 3.1200 0.4650 3.1800 0.5250 ;
        RECT 3.0150 0.1725 3.0750 0.2325 ;
        RECT 3.0150 0.8025 3.0750 0.8625 ;
        RECT 2.9100 0.3975 2.9700 0.4575 ;
        RECT 2.8050 0.1725 2.8650 0.2325 ;
        RECT 2.8050 0.7275 2.8650 0.7875 ;
        RECT 2.7000 0.4125 2.7600 0.4725 ;
        RECT 2.5950 0.1725 2.6550 0.2325 ;
        RECT 2.5950 0.8700 2.6550 0.9300 ;
        RECT 2.4900 0.4125 2.5500 0.4725 ;
        RECT 2.3850 0.7800 2.4450 0.8400 ;
        RECT 2.1750 0.2175 2.2350 0.2775 ;
        RECT 2.1750 0.8250 2.2350 0.8850 ;
        RECT 2.0700 0.5025 2.1300 0.5625 ;
        RECT 1.9650 0.2400 2.0250 0.3000 ;
        RECT 1.9650 0.7200 2.0250 0.7800 ;
        RECT 1.8600 0.5025 1.9200 0.5625 ;
        RECT 1.7550 0.2400 1.8150 0.3000 ;
        RECT 1.7550 0.7650 1.8150 0.8250 ;
        RECT 1.5450 0.1725 1.6050 0.2325 ;
        RECT 1.5450 0.7500 1.6050 0.8100 ;
        RECT 1.4400 0.4950 1.5000 0.5550 ;
        RECT 1.3350 0.1500 1.3950 0.2100 ;
        RECT 1.3350 0.8700 1.3950 0.9300 ;
        RECT 1.2300 0.4950 1.2900 0.5550 ;
        RECT 1.1250 0.1800 1.1850 0.2400 ;
        RECT 1.1250 0.7200 1.1850 0.7800 ;
        RECT 1.0200 0.4950 1.0800 0.5550 ;
        RECT 0.9150 0.1725 0.9750 0.2325 ;
        RECT 0.9150 0.8325 0.9750 0.8925 ;
        RECT 0.8100 0.3525 0.8700 0.4125 ;
        RECT 0.7050 0.1650 0.7650 0.2250 ;
        RECT 0.7050 0.8325 0.7650 0.8925 ;
        RECT 0.6000 0.6525 0.6600 0.7125 ;
        RECT 0.3900 0.6600 0.4500 0.7200 ;
        RECT 0.3825 0.4200 0.4425 0.4800 ;
        RECT 0.2850 0.1200 0.3450 0.1800 ;
        RECT 0.2850 0.8700 0.3450 0.9300 ;
        RECT 0.1875 0.4725 0.2475 0.5325 ;
        RECT 0.0750 0.2700 0.1350 0.3300 ;
        RECT 0.0750 0.8175 0.1350 0.8775 ;
        LAYER M1 ;
        RECT 6.0975 0.4350 6.2550 0.5550 ;
        RECT 6.1500 0.6525 6.2400 0.7875 ;
        RECT 5.9175 0.6525 6.1500 0.7275 ;
        RECT 5.9925 0.3675 6.0975 0.5550 ;
        RECT 5.9175 0.1650 6.0375 0.2700 ;
        RECT 5.8425 0.1650 5.9175 0.7275 ;
        RECT 5.6100 0.4575 5.8425 0.5550 ;
        RECT 5.7675 0.8025 5.8350 0.9000 ;
        RECT 5.6925 0.6375 5.7675 0.9000 ;
        RECT 5.2875 0.6375 5.6925 0.7125 ;
        RECT 5.1825 0.2625 5.6475 0.3375 ;
        RECT 5.1975 0.4125 5.5125 0.5550 ;
        RECT 5.2125 0.6375 5.2875 0.9000 ;
        RECT 5.0925 0.7950 5.2125 0.9000 ;
        RECT 5.1075 0.1950 5.1825 0.3375 ;
        RECT 4.4925 0.6450 5.1075 0.7200 ;
        RECT 4.7775 0.4650 5.0925 0.5700 ;
        RECT 4.8750 0.1500 5.0325 0.3600 ;
        RECT 4.6425 0.7950 4.9875 0.9000 ;
        RECT 4.4925 0.1500 4.7775 0.2550 ;
        RECT 4.5675 0.3300 4.7025 0.5700 ;
        RECT 4.4175 0.1500 4.4925 0.7200 ;
        RECT 4.1550 0.3225 4.4175 0.3975 ;
        RECT 4.1325 0.6450 4.4175 0.7200 ;
        RECT 4.0425 0.4800 4.3050 0.5700 ;
        RECT 4.1100 0.2775 4.1550 0.3975 ;
        RECT 4.0575 0.6450 4.1325 0.8250 ;
        RECT 4.0350 0.2775 4.1100 0.3900 ;
        RECT 3.9375 0.4650 4.0425 0.5700 ;
        RECT 3.7500 0.4425 3.8400 0.5400 ;
        RECT 3.1425 0.4425 3.7500 0.5325 ;
        RECT 3.6225 0.1950 3.7275 0.3675 ;
        RECT 3.6375 0.6075 3.7125 0.8700 ;
        RECT 3.2925 0.6075 3.6375 0.6975 ;
        RECT 3.3075 0.2775 3.6225 0.3675 ;
        RECT 3.2025 0.1950 3.3075 0.3675 ;
        RECT 3.2175 0.6075 3.2925 0.8700 ;
        RECT 3.0675 0.4425 3.1425 0.6450 ;
        RECT 2.6400 0.5550 3.0675 0.6450 ;
        RECT 2.8425 0.3750 2.9925 0.4800 ;
        RECT 2.7300 0.1500 2.9400 0.3000 ;
        RECT 2.4525 0.7200 2.8950 0.7950 ;
        RECT 2.4750 0.4050 2.8425 0.4800 ;
        RECT 2.4000 0.1875 2.4750 0.4800 ;
        RECT 2.3775 0.7200 2.4525 0.8925 ;
        RECT 2.1750 0.1875 2.4000 0.3075 ;
        RECT 2.1450 0.8175 2.3775 0.8925 ;
        RECT 2.0175 0.4800 2.3175 0.5850 ;
        RECT 2.0400 0.6600 2.2650 0.7425 ;
        RECT 1.9500 0.1650 2.1000 0.4050 ;
        RECT 1.9650 0.6600 2.0400 0.8250 ;
        RECT 1.8375 0.4800 1.9425 0.5850 ;
        RECT 1.7550 0.6600 1.8900 0.9000 ;
        RECT 1.7475 0.1500 1.8750 0.4050 ;
        RECT 1.5000 0.5100 1.8375 0.5850 ;
        RECT 1.5150 0.6675 1.6800 0.8700 ;
        RECT 1.5750 0.1500 1.6725 0.4050 ;
        RECT 1.5075 0.1500 1.5750 0.2550 ;
        RECT 1.4250 0.3300 1.5000 0.5850 ;
        RECT 1.3350 0.3300 1.4250 0.4125 ;
        RECT 1.2600 0.4875 1.3500 0.7575 ;
        RECT 1.1850 0.4875 1.2600 0.5925 ;
        RECT 1.0425 0.1500 1.2000 0.4125 ;
        RECT 1.1100 0.6675 1.1850 0.8100 ;
        RECT 1.0050 0.4875 1.1100 0.5925 ;
        RECT 0.6900 0.6675 1.1100 0.7425 ;
        RECT 0.8925 0.1500 1.0425 0.2550 ;
        RECT 0.5175 0.4875 1.0050 0.5625 ;
        RECT 0.5550 0.8175 1.0050 0.9000 ;
        RECT 0.6225 0.3300 0.9375 0.4125 ;
        RECT 0.7125 0.1500 0.8175 0.2550 ;
        RECT 0.4800 0.1500 0.7125 0.2325 ;
        RECT 0.5700 0.6375 0.6900 0.7425 ;
        RECT 0.5175 0.3075 0.6225 0.4125 ;
        RECT 0.4425 0.4875 0.5175 0.5775 ;
        RECT 0.1575 0.6600 0.4800 0.7650 ;
        RECT 0.3450 0.3900 0.4425 0.5775 ;
        RECT 0.1875 0.4425 0.3450 0.5775 ;
        RECT 0.1125 0.2625 0.2850 0.3375 ;
        RECT 0.1125 0.6600 0.1575 0.9000 ;
        RECT 0.0375 0.2625 0.1125 0.9000 ;
        LAYER VIA1 ;
        RECT 5.8425 0.6075 5.9175 0.6825 ;
        RECT 4.9500 0.4950 5.0250 0.5700 ;
        RECT 4.9125 0.1650 4.9875 0.2400 ;
        RECT 4.7625 0.8100 4.8375 0.8850 ;
        RECT 2.8800 0.3900 2.9550 0.4650 ;
        RECT 2.7900 0.1650 2.8650 0.2400 ;
        RECT 2.6850 0.5625 2.7600 0.6375 ;
        RECT 2.1750 0.4950 2.2500 0.5700 ;
        RECT 2.0175 0.6600 2.0925 0.7350 ;
        RECT 1.9875 0.3150 2.0625 0.3900 ;
        RECT 1.7850 0.7950 1.8600 0.8700 ;
        RECT 1.7700 0.2100 1.8450 0.2850 ;
        RECT 1.5750 0.2850 1.6500 0.3600 ;
        RECT 1.5600 0.6750 1.6350 0.7500 ;
        RECT 1.3800 0.3375 1.4550 0.4125 ;
        RECT 1.0875 0.3225 1.1625 0.3975 ;
        RECT 1.0425 0.6675 1.1175 0.7425 ;
        RECT 0.8250 0.8175 0.9000 0.8925 ;
        RECT 0.6975 0.1575 0.7725 0.2325 ;
        RECT 0.5625 0.3375 0.6375 0.4125 ;
        RECT 0.1650 0.2625 0.2400 0.3375 ;
        LAYER M2 ;
        RECT 5.8275 0.5625 5.9325 0.7200 ;
        RECT 5.1000 0.5625 5.8275 0.6375 ;
        RECT 5.0250 0.4950 5.1000 0.6375 ;
        RECT 4.5525 0.1650 5.0325 0.2400 ;
        RECT 4.8975 0.4950 5.0250 0.5700 ;
        RECT 4.5525 0.8100 4.8825 0.8850 ;
        RECT 4.4775 0.1650 4.5525 0.8850 ;
        RECT 2.9925 0.8100 4.4775 0.8850 ;
        RECT 2.9175 0.3750 2.9925 0.8850 ;
        RECT 2.8425 0.3750 2.9175 0.4800 ;
        RECT 1.8975 0.8100 2.9175 0.8850 ;
        RECT 1.8525 0.1650 2.9100 0.2400 ;
        RECT 2.6850 0.3150 2.7600 0.7350 ;
        RECT 2.0400 0.3150 2.6850 0.3900 ;
        RECT 1.9725 0.6600 2.6850 0.7350 ;
        RECT 1.6500 0.4950 2.2950 0.5700 ;
        RECT 1.9350 0.3150 2.0400 0.4200 ;
        RECT 1.7475 0.7800 1.8975 0.8850 ;
        RECT 1.7475 0.1650 1.8525 0.3300 ;
        RECT 1.5750 0.2400 1.6500 0.7875 ;
        RECT 1.5450 0.6375 1.5750 0.7875 ;
        RECT 1.4175 0.3075 1.5000 0.4125 ;
        RECT 1.3350 0.1575 1.4175 0.4125 ;
        RECT 0.9525 0.1575 1.3350 0.2325 ;
        RECT 1.1325 0.3150 1.2075 0.4200 ;
        RECT 1.0275 0.3150 1.1325 0.7875 ;
        RECT 0.8775 0.1575 0.9525 0.9000 ;
        RECT 0.6525 0.1575 0.8775 0.2325 ;
        RECT 0.7800 0.7950 0.8775 0.9000 ;
        RECT 0.5100 0.3375 0.6825 0.4125 ;
        RECT 0.4350 0.2625 0.5100 0.4125 ;
        RECT 0.1200 0.2625 0.4350 0.3375 ;
    END
END XNR4_0111


MACRO XOR2_0011
    CLASS CORE ;
    FOREIGN XOR2_0011 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.8900 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 1.7775 0.3075 1.8525 0.7500 ;
        RECT 1.6125 0.3075 1.7775 0.3825 ;
        RECT 1.6125 0.6750 1.7775 0.7500 ;
        RECT 1.5375 0.2175 1.6125 0.3825 ;
        RECT 1.5375 0.6750 1.6125 0.8175 ;
        END
    END Z
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.0950 0.4125 1.5300 0.4875 ;
        RECT 1.0200 0.3750 1.0950 0.4875 ;
        VIA 1.2600 0.4500 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.1350 0.4125 0.6000 0.4875 ;
        VIA 0.3150 0.4500 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.8450 -0.0750 1.8900 0.0750 ;
        RECT 1.7250 -0.0750 1.8450 0.2250 ;
        RECT 1.4025 -0.0750 1.7250 0.0750 ;
        RECT 1.2975 -0.0750 1.4025 0.2550 ;
        RECT 0.3600 -0.0750 1.2975 0.0750 ;
        RECT 0.2700 -0.0750 0.3600 0.2250 ;
        RECT 0.0000 -0.0750 0.2700 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.8450 0.9750 1.8900 1.1250 ;
        RECT 1.7250 0.8250 1.8450 1.1250 ;
        RECT 1.4250 0.9750 1.7250 1.1250 ;
        RECT 1.3050 0.8700 1.4250 1.1250 ;
        RECT 0.3750 0.9750 1.3050 1.1250 ;
        RECT 0.2550 0.8175 0.3750 1.1250 ;
        RECT 0.0000 0.9750 0.2550 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.7550 0.1575 1.8150 0.2175 ;
        RECT 1.7550 0.8325 1.8150 0.8925 ;
        RECT 1.6425 0.4950 1.7025 0.5550 ;
        RECT 1.5450 0.2925 1.6050 0.3525 ;
        RECT 1.5450 0.7200 1.6050 0.7800 ;
        RECT 1.4400 0.4950 1.5000 0.5550 ;
        RECT 1.3350 0.1650 1.3950 0.2250 ;
        RECT 1.3350 0.8700 1.3950 0.9300 ;
        RECT 1.2300 0.4650 1.2900 0.5250 ;
        RECT 1.1250 0.1800 1.1850 0.2400 ;
        RECT 1.1250 0.7275 1.1850 0.7875 ;
        RECT 1.0125 0.4650 1.0725 0.5250 ;
        RECT 0.9150 0.1800 0.9750 0.2400 ;
        RECT 0.9150 0.8325 0.9750 0.8925 ;
        RECT 0.8100 0.5025 0.8700 0.5625 ;
        RECT 0.7050 0.1800 0.7650 0.2400 ;
        RECT 0.7050 0.8325 0.7650 0.8925 ;
        RECT 0.6000 0.6525 0.6600 0.7125 ;
        RECT 0.3900 0.3450 0.4500 0.4050 ;
        RECT 0.3900 0.6600 0.4500 0.7200 ;
        RECT 0.2850 0.1350 0.3450 0.1950 ;
        RECT 0.2850 0.8400 0.3450 0.9000 ;
        RECT 0.1875 0.4800 0.2475 0.5400 ;
        RECT 0.0750 0.1800 0.1350 0.2400 ;
        RECT 0.0750 0.8175 0.1350 0.8775 ;
        LAYER M1 ;
        RECT 1.4625 0.4650 1.7025 0.5850 ;
        RECT 1.3725 0.4650 1.4625 0.7950 ;
        RECT 1.2600 0.6300 1.3725 0.7950 ;
        RECT 1.1475 0.3300 1.2975 0.5550 ;
        RECT 0.8775 0.1500 1.2225 0.2550 ;
        RECT 1.1100 0.6600 1.1850 0.8250 ;
        RECT 0.6825 0.6600 1.1100 0.7350 ;
        RECT 0.9975 0.3300 1.0725 0.5550 ;
        RECT 0.6300 0.8100 1.0050 0.9000 ;
        RECT 0.3525 0.3300 0.9975 0.4050 ;
        RECT 0.7725 0.4800 0.8925 0.5850 ;
        RECT 0.4950 0.1500 0.7950 0.2550 ;
        RECT 0.5025 0.4800 0.7725 0.5550 ;
        RECT 0.5775 0.6300 0.6825 0.7350 ;
        RECT 0.4275 0.4800 0.5025 0.7350 ;
        RECT 0.1575 0.6600 0.4275 0.7350 ;
        RECT 0.2775 0.3300 0.3525 0.5700 ;
        RECT 0.1875 0.4500 0.2775 0.5700 ;
        RECT 0.1125 0.6600 0.1575 0.9000 ;
        RECT 0.1125 0.1500 0.1425 0.2700 ;
        RECT 0.0375 0.1500 0.1125 0.9000 ;
        LAYER VIA1 ;
        RECT 1.2600 0.6750 1.3350 0.7500 ;
        RECT 0.9450 0.6600 1.0200 0.7350 ;
        RECT 0.9225 0.1650 0.9975 0.2400 ;
        RECT 0.7650 0.8100 0.8400 0.8850 ;
        RECT 0.6825 0.1650 0.7575 0.2400 ;
        LAYER M2 ;
        RECT 1.2600 0.6300 1.3350 0.8850 ;
        RECT 0.7950 0.8100 1.2600 0.8850 ;
        RECT 0.9450 0.6600 1.0650 0.7350 ;
        RECT 0.9450 0.1500 1.0425 0.2550 ;
        RECT 0.8700 0.1500 0.9450 0.7350 ;
        RECT 0.7200 0.1500 0.7950 0.8850 ;
        RECT 0.6450 0.1500 0.7200 0.2550 ;
    END
END XOR2_0011


MACRO XOR2_0111
    CLASS CORE ;
    FOREIGN XOR2_0111 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.3600 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 2.6775 0.2400 2.9925 0.7500 ;
        VIA 2.8350 0.3225 VIA12_slot ;
        VIA 2.8350 0.6675 VIA12_slot ;
        END
    END Z
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 2.0775 0.4425 2.1525 0.6375 ;
        RECT 1.6125 0.5625 2.0775 0.6375 ;
        VIA 2.1150 0.5250 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.6275 0.4125 1.7775 0.4875 ;
        RECT 1.5525 0.3225 1.6275 0.4875 ;
        RECT 1.0950 0.3225 1.5525 0.4050 ;
        RECT 1.0200 0.3225 1.0950 0.4875 ;
        RECT 0.4725 0.4125 1.0200 0.4875 ;
        RECT 0.3675 0.2625 0.4725 0.4875 ;
        VIA 1.6650 0.4500 VIA12_square ;
        VIA 0.9525 0.4500 VIA12_square ;
        VIA 0.4200 0.3375 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 3.2925 -0.0750 3.3600 0.0750 ;
        RECT 3.2175 -0.0750 3.2925 0.3150 ;
        RECT 2.8950 -0.0750 3.2175 0.0750 ;
        RECT 2.7750 -0.0750 2.8950 0.1950 ;
        RECT 2.4525 -0.0750 2.7750 0.0750 ;
        RECT 2.3775 -0.0750 2.4525 0.3075 ;
        RECT 2.0625 -0.0750 2.3775 0.0750 ;
        RECT 1.9575 -0.0750 2.0625 0.2475 ;
        RECT 1.0050 -0.0750 1.9575 0.0750 ;
        RECT 0.8850 -0.0750 1.0050 0.1875 ;
        RECT 0.3750 -0.0750 0.8850 0.0750 ;
        RECT 0.2550 -0.0750 0.3750 0.2250 ;
        RECT 0.0000 -0.0750 0.2550 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 3.2925 0.9750 3.3600 1.1250 ;
        RECT 3.2175 0.6375 3.2925 1.1250 ;
        RECT 2.8875 0.9750 3.2175 1.1250 ;
        RECT 2.7825 0.8025 2.8875 1.1250 ;
        RECT 2.4750 0.9750 2.7825 1.1250 ;
        RECT 2.3550 0.6600 2.4750 1.1250 ;
        RECT 2.0550 0.9750 2.3550 1.1250 ;
        RECT 1.9350 0.8025 2.0550 1.1250 ;
        RECT 0.7875 0.9750 1.9350 1.1250 ;
        RECT 0.6825 0.7875 0.7875 1.1250 ;
        RECT 0.3675 0.9750 0.6825 1.1250 ;
        RECT 0.2625 0.8100 0.3675 1.1250 ;
        RECT 0.0000 0.9750 0.2625 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 3.2250 0.2250 3.2850 0.2850 ;
        RECT 3.2250 0.6675 3.2850 0.7275 ;
        RECT 3.2250 0.8325 3.2850 0.8925 ;
        RECT 3.1200 0.4650 3.1800 0.5250 ;
        RECT 3.0150 0.2250 3.0750 0.2850 ;
        RECT 3.0150 0.7575 3.0750 0.8175 ;
        RECT 2.9100 0.4650 2.9700 0.5250 ;
        RECT 2.8050 0.1275 2.8650 0.1875 ;
        RECT 2.8050 0.8325 2.8650 0.8925 ;
        RECT 2.7000 0.4650 2.7600 0.5250 ;
        RECT 2.5950 0.2250 2.6550 0.2850 ;
        RECT 2.5950 0.7575 2.6550 0.8175 ;
        RECT 2.4900 0.4650 2.5500 0.5250 ;
        RECT 2.3850 0.2175 2.4450 0.2775 ;
        RECT 2.3850 0.6675 2.4450 0.7275 ;
        RECT 2.3850 0.8325 2.4450 0.8925 ;
        RECT 2.2800 0.4875 2.3400 0.5475 ;
        RECT 2.1750 0.3075 2.2350 0.3675 ;
        RECT 2.1750 0.7275 2.2350 0.7875 ;
        RECT 2.0700 0.4875 2.1300 0.5475 ;
        RECT 1.9650 0.1575 2.0250 0.2175 ;
        RECT 1.9650 0.8100 2.0250 0.8700 ;
        RECT 1.7550 0.6525 1.8150 0.7125 ;
        RECT 1.6500 0.4500 1.7100 0.5100 ;
        RECT 1.5450 0.1725 1.6050 0.2325 ;
        RECT 1.5450 0.8250 1.6050 0.8850 ;
        RECT 1.4400 0.4875 1.5000 0.5475 ;
        RECT 1.3350 0.2325 1.3950 0.2925 ;
        RECT 1.3350 0.8175 1.3950 0.8775 ;
        RECT 1.2300 0.6450 1.2900 0.7050 ;
        RECT 1.1250 0.2400 1.1850 0.3000 ;
        RECT 1.1250 0.8175 1.1850 0.8775 ;
        RECT 1.0200 0.4650 1.0800 0.5250 ;
        RECT 0.9150 0.1275 0.9750 0.1875 ;
        RECT 0.8100 0.4650 0.8700 0.5250 ;
        RECT 0.7050 0.2700 0.7650 0.3300 ;
        RECT 0.7050 0.8175 0.7650 0.8775 ;
        RECT 0.6000 0.4800 0.6600 0.5400 ;
        RECT 0.4950 0.8175 0.5550 0.8775 ;
        RECT 0.3900 0.4800 0.4500 0.5400 ;
        RECT 0.2850 0.1575 0.3450 0.2175 ;
        RECT 0.2850 0.8325 0.3450 0.8925 ;
        RECT 0.1875 0.4725 0.2475 0.5325 ;
        RECT 0.0750 0.2100 0.1350 0.2700 ;
        RECT 0.0750 0.7350 0.1350 0.7950 ;
        LAYER M1 ;
        RECT 2.4375 0.4425 3.2100 0.5475 ;
        RECT 2.9925 0.1950 3.0975 0.3675 ;
        RECT 3.0075 0.6225 3.0825 0.8700 ;
        RECT 2.6625 0.6225 3.0075 0.7125 ;
        RECT 2.6775 0.2775 2.9925 0.3675 ;
        RECT 2.5725 0.1950 2.6775 0.3675 ;
        RECT 2.5875 0.6225 2.6625 0.8700 ;
        RECT 2.2575 0.4650 2.3625 0.5700 ;
        RECT 2.1900 0.2775 2.2650 0.3900 ;
        RECT 1.9950 0.4800 2.2575 0.5700 ;
        RECT 2.1675 0.6450 2.2425 0.8250 ;
        RECT 2.1450 0.2775 2.1900 0.3975 ;
        RECT 1.8825 0.6450 2.1675 0.7200 ;
        RECT 1.8825 0.3225 2.1450 0.3975 ;
        RECT 1.8075 0.1500 1.8825 0.7200 ;
        RECT 1.5225 0.1500 1.8075 0.2550 ;
        RECT 1.1925 0.6450 1.8075 0.7200 ;
        RECT 1.5975 0.3300 1.7325 0.5700 ;
        RECT 1.3125 0.7950 1.6575 0.9000 ;
        RECT 1.2075 0.4650 1.5225 0.5700 ;
        RECT 1.2675 0.1500 1.4250 0.3600 ;
        RECT 1.0875 0.7950 1.2075 0.9000 ;
        RECT 1.1175 0.1950 1.1925 0.3375 ;
        RECT 0.6600 0.2625 1.1175 0.3375 ;
        RECT 1.0125 0.6375 1.0875 0.9000 ;
        RECT 0.8100 0.4125 1.0800 0.5550 ;
        RECT 0.6075 0.6375 1.0125 0.7125 ;
        RECT 0.4575 0.4500 0.6900 0.5550 ;
        RECT 0.5325 0.6375 0.6075 0.9000 ;
        RECT 0.4725 0.7950 0.5325 0.9000 ;
        RECT 0.3075 0.3000 0.5025 0.3750 ;
        RECT 0.3825 0.4500 0.4575 0.7200 ;
        RECT 0.1350 0.6450 0.3825 0.7200 ;
        RECT 0.2325 0.3000 0.3075 0.5625 ;
        RECT 0.1875 0.4425 0.2325 0.5625 ;
        RECT 0.1125 0.1800 0.1425 0.3000 ;
        RECT 0.1125 0.6450 0.1350 0.8325 ;
        RECT 0.0375 0.1800 0.1125 0.8325 ;
        LAYER VIA1 ;
        RECT 2.4750 0.4575 2.5500 0.5325 ;
        RECT 1.4625 0.8100 1.5375 0.8850 ;
        RECT 1.3125 0.1650 1.3875 0.2400 ;
        RECT 1.2750 0.4950 1.3500 0.5700 ;
        RECT 0.3825 0.5625 0.4575 0.6375 ;
        LAYER M2 ;
        RECT 2.3325 0.4200 2.5650 0.5700 ;
        RECT 2.2575 0.1650 2.3325 0.8850 ;
        RECT 1.2675 0.1650 2.2575 0.2400 ;
        RECT 1.4175 0.8100 2.2575 0.8850 ;
        RECT 1.2600 0.4950 1.4025 0.5700 ;
        RECT 1.1850 0.4950 1.2600 0.6375 ;
        RECT 0.3075 0.5625 1.1850 0.6375 ;
    END
END XOR2_0111


MACRO XOR2_1000
    CLASS CORE ;
    FOREIGN XOR2_1000 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.5100 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 5.8800 0.3150 6.0375 0.4350 ;
        RECT 5.8800 0.6150 6.0375 0.7350 ;
        RECT 5.5650 0.3150 5.8800 0.7350 ;
        RECT 5.4075 0.3150 5.5650 0.4350 ;
        RECT 5.4075 0.6150 5.5650 0.7350 ;
        VIA 5.8800 0.3750 VIA12_slot ;
        VIA 5.8800 0.6750 VIA12_slot ;
        VIA 5.5650 0.3750 VIA12_slot ;
        VIA 5.5650 0.6750 VIA12_slot ;
        END
    END Z
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.1100 0.4350 1.2225 0.6375 ;
        RECT 0.6000 0.5625 1.1100 0.6375 ;
        VIA 1.1700 0.5175 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 3.2325 0.4125 3.9975 0.4875 ;
        RECT 3.1275 0.4125 3.2325 0.6075 ;
        VIA 3.8775 0.4500 VIA12_square ;
        VIA 3.1800 0.5175 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 3.5400 -0.0750 6.5100 0.0750 ;
        RECT 3.3900 -0.0750 3.5400 0.2175 ;
        RECT 3.1050 -0.0750 3.3900 0.0750 ;
        RECT 2.9850 -0.0750 3.1050 0.2250 ;
        RECT 2.6850 -0.0750 2.9850 0.0750 ;
        RECT 2.5650 -0.0750 2.6850 0.2325 ;
        RECT 2.2650 -0.0750 2.5650 0.0750 ;
        RECT 2.1450 -0.0750 2.2650 0.2325 ;
        RECT 1.8450 -0.0750 2.1450 0.0750 ;
        RECT 1.7250 -0.0750 1.8450 0.2325 ;
        RECT 1.4250 -0.0750 1.7250 0.0750 ;
        RECT 1.3050 -0.0750 1.4250 0.2325 ;
        RECT 1.0050 -0.0750 1.3050 0.0750 ;
        RECT 0.8850 -0.0750 1.0050 0.2325 ;
        RECT 0.5775 -0.0750 0.8850 0.0750 ;
        RECT 0.4725 -0.0750 0.5775 0.2325 ;
        RECT 0.1650 -0.0750 0.4725 0.0750 ;
        RECT 0.0450 -0.0750 0.1650 0.2325 ;
        RECT 0.0000 -0.0750 0.0450 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 3.5250 0.9750 6.5100 1.1250 ;
        RECT 3.4050 0.8325 3.5250 1.1250 ;
        RECT 3.1200 0.9750 3.4050 1.1250 ;
        RECT 2.9700 0.8325 3.1200 1.1250 ;
        RECT 2.6850 0.9750 2.9700 1.1250 ;
        RECT 2.5650 0.8400 2.6850 1.1250 ;
        RECT 2.2650 0.9750 2.5650 1.1250 ;
        RECT 2.1450 0.8400 2.2650 1.1250 ;
        RECT 1.8450 0.9750 2.1450 1.1250 ;
        RECT 1.7250 0.8400 1.8450 1.1250 ;
        RECT 1.4250 0.9750 1.7250 1.1250 ;
        RECT 1.3050 0.8400 1.4250 1.1250 ;
        RECT 1.0050 0.9750 1.3050 1.1250 ;
        RECT 0.8850 0.8400 1.0050 1.1250 ;
        RECT 0.5850 0.9750 0.8850 1.1250 ;
        RECT 0.4650 0.8400 0.5850 1.1250 ;
        RECT 0.1650 0.9750 0.4650 1.1250 ;
        RECT 0.0450 0.8100 0.1650 1.1250 ;
        RECT 0.0000 0.9750 0.0450 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 6.3750 0.3075 6.4350 0.3675 ;
        RECT 6.3750 0.6750 6.4350 0.7350 ;
        RECT 6.2700 0.4950 6.3300 0.5550 ;
        RECT 6.1650 0.1575 6.2250 0.2175 ;
        RECT 6.1650 0.8325 6.2250 0.8925 ;
        RECT 6.0600 0.4950 6.1200 0.5550 ;
        RECT 5.9550 0.3225 6.0150 0.3825 ;
        RECT 5.9550 0.6750 6.0150 0.7350 ;
        RECT 5.8500 0.4950 5.9100 0.5550 ;
        RECT 5.7450 0.1575 5.8050 0.2175 ;
        RECT 5.7450 0.8325 5.8050 0.8925 ;
        RECT 5.6400 0.4950 5.7000 0.5550 ;
        RECT 5.5350 0.3225 5.5950 0.3825 ;
        RECT 5.5350 0.6750 5.5950 0.7350 ;
        RECT 5.4300 0.4950 5.4900 0.5550 ;
        RECT 5.3250 0.1575 5.3850 0.2175 ;
        RECT 5.3250 0.8325 5.3850 0.8925 ;
        RECT 5.2200 0.4950 5.2800 0.5550 ;
        RECT 5.1150 0.2625 5.1750 0.3225 ;
        RECT 5.1150 0.6750 5.1750 0.7350 ;
        RECT 5.0100 0.4800 5.0700 0.5400 ;
        RECT 4.9050 0.3000 4.9650 0.3600 ;
        RECT 4.9050 0.6675 4.9650 0.7275 ;
        RECT 4.8000 0.4800 4.8600 0.5400 ;
        RECT 4.6950 0.1575 4.7550 0.2175 ;
        RECT 4.6950 0.8325 4.7550 0.8925 ;
        RECT 4.5900 0.4800 4.6500 0.5400 ;
        RECT 4.4850 0.3000 4.5450 0.3600 ;
        RECT 4.4850 0.6675 4.5450 0.7275 ;
        RECT 4.3800 0.4800 4.4400 0.5400 ;
        RECT 4.2750 0.1575 4.3350 0.2175 ;
        RECT 4.2750 0.8325 4.3350 0.8925 ;
        RECT 4.1700 0.4800 4.2300 0.5400 ;
        RECT 4.0650 0.3000 4.1250 0.3600 ;
        RECT 4.0650 0.6825 4.1250 0.7425 ;
        RECT 3.9600 0.4800 4.0200 0.5400 ;
        RECT 3.8550 0.1875 3.9150 0.2475 ;
        RECT 3.8550 0.8025 3.9150 0.8625 ;
        RECT 3.6450 0.3075 3.7050 0.3675 ;
        RECT 3.6450 0.6900 3.7050 0.7500 ;
        RECT 3.5400 0.4875 3.6000 0.5475 ;
        RECT 3.4350 0.1575 3.4950 0.2175 ;
        RECT 3.4350 0.8325 3.4950 0.8925 ;
        RECT 3.3300 0.4875 3.3900 0.5475 ;
        RECT 3.2250 0.3075 3.2850 0.3675 ;
        RECT 3.2250 0.6900 3.2850 0.7500 ;
        RECT 3.1200 0.4875 3.1800 0.5475 ;
        RECT 3.0150 0.1425 3.0750 0.2025 ;
        RECT 3.0150 0.8325 3.0750 0.8925 ;
        RECT 2.9100 0.4875 2.9700 0.5475 ;
        RECT 2.8050 0.2925 2.8650 0.3525 ;
        RECT 2.8050 0.7200 2.8650 0.7800 ;
        RECT 2.7000 0.4875 2.7600 0.5475 ;
        RECT 2.5950 0.1650 2.6550 0.2250 ;
        RECT 2.5950 0.8475 2.6550 0.9075 ;
        RECT 2.4900 0.4875 2.5500 0.5475 ;
        RECT 2.3850 0.3075 2.4450 0.3675 ;
        RECT 2.3850 0.6825 2.4450 0.7425 ;
        RECT 2.2800 0.4875 2.3400 0.5475 ;
        RECT 2.1750 0.1650 2.2350 0.2250 ;
        RECT 2.1750 0.8475 2.2350 0.9075 ;
        RECT 2.0700 0.4875 2.1300 0.5475 ;
        RECT 1.9650 0.2925 2.0250 0.3525 ;
        RECT 1.9650 0.7350 2.0250 0.7950 ;
        RECT 1.8600 0.4875 1.9200 0.5475 ;
        RECT 1.7550 0.1650 1.8150 0.2250 ;
        RECT 1.7550 0.8475 1.8150 0.9075 ;
        RECT 1.6500 0.4875 1.7100 0.5475 ;
        RECT 1.5450 0.3075 1.6050 0.3675 ;
        RECT 1.5450 0.6900 1.6050 0.7500 ;
        RECT 1.4400 0.4875 1.5000 0.5475 ;
        RECT 1.3350 0.1650 1.3950 0.2250 ;
        RECT 1.3350 0.8475 1.3950 0.9075 ;
        RECT 1.2300 0.4875 1.2900 0.5475 ;
        RECT 1.1250 0.3075 1.1850 0.3675 ;
        RECT 1.1250 0.6900 1.1850 0.7500 ;
        RECT 1.0200 0.4875 1.0800 0.5475 ;
        RECT 0.9150 0.1650 0.9750 0.2250 ;
        RECT 0.9150 0.8475 0.9750 0.9075 ;
        RECT 0.8100 0.4875 0.8700 0.5475 ;
        RECT 0.7050 0.3075 0.7650 0.3675 ;
        RECT 0.7050 0.6900 0.7650 0.7500 ;
        RECT 0.6000 0.4875 0.6600 0.5475 ;
        RECT 0.4950 0.1500 0.5550 0.2100 ;
        RECT 0.4950 0.8475 0.5550 0.9075 ;
        RECT 0.3900 0.4875 0.4500 0.5475 ;
        RECT 0.2850 0.2925 0.3450 0.3525 ;
        RECT 0.2850 0.7350 0.3450 0.7950 ;
        RECT 0.1800 0.4875 0.2400 0.5475 ;
        RECT 0.0750 0.1650 0.1350 0.2250 ;
        RECT 0.0750 0.8175 0.1350 0.8775 ;
        LAYER M1 ;
        RECT 6.3450 0.2775 6.4650 0.4125 ;
        RECT 6.3600 0.6375 6.4425 0.7875 ;
        RECT 5.3400 0.4875 6.3900 0.5625 ;
        RECT 5.4075 0.6375 6.3600 0.7350 ;
        RECT 5.4075 0.3075 6.3450 0.4125 ;
        RECT 5.4525 0.1500 6.2775 0.2250 ;
        RECT 5.4075 0.8250 6.2550 0.9000 ;
        RECT 5.2875 0.1500 5.4525 0.2325 ;
        RECT 5.1825 0.3075 5.4075 0.3825 ;
        RECT 5.1375 0.6600 5.4075 0.7350 ;
        RECT 5.2425 0.8175 5.4075 0.9000 ;
        RECT 5.1450 0.4575 5.3400 0.5850 ;
        RECT 5.1075 0.1500 5.1825 0.3825 ;
        RECT 5.0625 0.6600 5.1375 0.9000 ;
        RECT 3.9300 0.1500 5.1075 0.2250 ;
        RECT 4.9650 0.4500 5.0700 0.5700 ;
        RECT 3.9225 0.8250 5.0625 0.9000 ;
        RECT 4.0350 0.3000 4.9950 0.3750 ;
        RECT 4.4025 0.6450 4.9875 0.7500 ;
        RECT 3.9300 0.4500 4.9650 0.5400 ;
        RECT 4.0350 0.6750 4.4025 0.7500 ;
        RECT 3.8250 0.1500 3.9300 0.2850 ;
        RECT 3.8250 0.3750 3.9300 0.5400 ;
        RECT 3.8475 0.7575 3.9225 0.9000 ;
        RECT 3.6750 0.3075 3.7500 0.7575 ;
        RECT 3.1875 0.3075 3.6750 0.3825 ;
        RECT 3.1875 0.6525 3.6750 0.7575 ;
        RECT 3.0825 0.4575 3.6000 0.5775 ;
        RECT 2.8425 0.4725 3.0000 0.5775 ;
        RECT 2.7975 0.2625 2.8725 0.3825 ;
        RECT 2.7975 0.6675 2.8725 0.8325 ;
        RECT 1.8600 0.4575 2.8425 0.5775 ;
        RECT 2.0325 0.3075 2.7975 0.3825 ;
        RECT 2.0325 0.6675 2.7975 0.7425 ;
        RECT 1.9575 0.2250 2.0325 0.3825 ;
        RECT 1.9575 0.6675 2.0325 0.8400 ;
        RECT 1.7850 0.3075 1.8600 0.7575 ;
        RECT 0.3525 0.3075 1.7850 0.3825 ;
        RECT 0.3525 0.6825 1.7850 0.7575 ;
        RECT 0.1500 0.4575 1.7100 0.5775 ;
        RECT 0.2775 0.2325 0.3525 0.3825 ;
        RECT 0.2775 0.6825 0.3525 0.8400 ;
        LAYER VIA1 ;
        RECT 5.3325 0.1575 5.4075 0.2325 ;
        RECT 5.2875 0.8175 5.3625 0.8925 ;
        RECT 5.1825 0.4800 5.2575 0.5550 ;
        RECT 4.4475 0.6675 4.5225 0.7425 ;
        RECT 4.2225 0.3000 4.2975 0.3750 ;
        RECT 3.6750 0.5625 3.7500 0.6375 ;
        RECT 2.8575 0.4800 2.9325 0.5550 ;
        RECT 2.7975 0.7125 2.8725 0.7875 ;
        RECT 2.6400 0.3075 2.7150 0.3825 ;
        RECT 2.4300 0.4875 2.5050 0.5625 ;
        LAYER M2 ;
        RECT 5.9100 0.3150 6.0375 0.4350 ;
        RECT 5.9100 0.6150 6.0375 0.7350 ;
        RECT 5.4075 0.3150 5.5350 0.4350 ;
        RECT 5.4075 0.6150 5.5350 0.7350 ;
        RECT 5.2875 0.1125 5.4525 0.2325 ;
        RECT 5.2425 0.8175 5.4075 0.9375 ;
        RECT 2.7150 0.1125 5.2875 0.1875 ;
        RECT 5.1825 0.4275 5.2575 0.6225 ;
        RECT 2.5050 0.8625 5.2425 0.9375 ;
        RECT 4.5375 0.4275 5.1825 0.5025 ;
        RECT 4.4325 0.6225 4.5450 0.7875 ;
        RECT 4.4625 0.4275 4.5375 0.5475 ;
        RECT 4.3575 0.4725 4.4625 0.5475 ;
        RECT 2.7150 0.7125 4.4325 0.7875 ;
        RECT 4.2825 0.4725 4.3575 0.6375 ;
        RECT 4.1775 0.2625 4.3425 0.3900 ;
        RECT 3.6150 0.5625 4.2825 0.6375 ;
        RECT 2.9475 0.2625 4.1775 0.3375 ;
        RECT 2.8425 0.2625 2.9475 0.6000 ;
        RECT 2.6400 0.1125 2.7150 0.7875 ;
        RECT 2.4300 0.3825 2.5050 0.9375 ;
    END
END XOR2_1000


MACRO XOR2_1010
    CLASS CORE ;
    FOREIGN XOR2_1010 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.4700 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 0.7875 0.8625 1.2525 0.9375 ;
        RECT 0.7125 0.1650 0.7875 0.9375 ;
        RECT 0.5925 0.1650 0.7125 0.2400 ;
        VIA 0.7500 0.8475 VIA12_square ;
        VIA 0.6750 0.2025 VIA12_square ;
        END
    END Z
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.3125 0.3675 1.4175 0.6825 ;
        RECT 1.2300 0.3675 1.3125 0.5550 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.1275 0.5625 0.5925 0.6375 ;
        VIA 0.3150 0.6000 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.4250 -0.0750 1.4700 0.0750 ;
        RECT 1.3050 -0.0750 1.4250 0.2550 ;
        RECT 0.3750 -0.0750 1.3050 0.0750 ;
        RECT 0.2550 -0.0750 0.3750 0.2400 ;
        RECT 0.0000 -0.0750 0.2550 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 1.4250 0.9750 1.4700 1.1250 ;
        RECT 1.3050 0.7575 1.4250 1.1250 ;
        RECT 0.3750 0.9750 1.3050 1.1250 ;
        RECT 0.2550 0.8625 0.3750 1.1250 ;
        RECT 0.0000 0.9750 0.2550 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 1.3350 0.1650 1.3950 0.2250 ;
        RECT 1.3350 0.7875 1.3950 0.8475 ;
        RECT 1.2300 0.4650 1.2900 0.5250 ;
        RECT 1.1250 0.1800 1.1850 0.2400 ;
        RECT 1.1250 0.7275 1.1850 0.7875 ;
        RECT 1.0200 0.4500 1.0800 0.5100 ;
        RECT 0.9150 0.1800 0.9750 0.2400 ;
        RECT 0.9150 0.8325 0.9750 0.8925 ;
        RECT 0.8100 0.5025 0.8700 0.5625 ;
        RECT 0.7050 0.1800 0.7650 0.2400 ;
        RECT 0.7050 0.8325 0.7650 0.8925 ;
        RECT 0.6000 0.6600 0.6600 0.7200 ;
        RECT 0.3900 0.3450 0.4500 0.4050 ;
        RECT 0.3900 0.6600 0.4500 0.7200 ;
        RECT 0.2850 0.1500 0.3450 0.2100 ;
        RECT 0.2850 0.8700 0.3450 0.9300 ;
        RECT 0.1875 0.5250 0.2475 0.5850 ;
        RECT 0.0750 0.1875 0.1350 0.2475 ;
        RECT 0.0750 0.8175 0.1350 0.8775 ;
        LAYER M1 ;
        RECT 0.8700 0.1500 1.2150 0.2550 ;
        RECT 1.1175 0.6600 1.1925 0.8250 ;
        RECT 0.5625 0.6600 1.1175 0.7350 ;
        RECT 1.0125 0.3375 1.0875 0.5400 ;
        RECT 0.1425 0.3375 1.0125 0.4125 ;
        RECT 0.6000 0.8100 1.0050 0.9000 ;
        RECT 0.4575 0.4950 0.9000 0.5700 ;
        RECT 0.4650 0.1500 0.7950 0.2550 ;
        RECT 0.3525 0.4950 0.4575 0.7650 ;
        RECT 0.1875 0.4950 0.3525 0.6375 ;
        RECT 0.1125 0.7950 0.1575 0.9000 ;
        RECT 0.1125 0.1575 0.1425 0.4125 ;
        RECT 0.0375 0.1575 0.1125 0.9000 ;
        LAYER VIA1 ;
        RECT 0.9075 0.1650 0.9825 0.2400 ;
        RECT 0.9075 0.6600 0.9825 0.7350 ;
        LAYER M2 ;
        RECT 0.9675 0.1275 0.9975 0.2775 ;
        RECT 0.9675 0.6225 0.9975 0.7725 ;
        RECT 0.8925 0.1275 0.9675 0.7725 ;
    END
END XOR2_1010


MACRO XOR3_0011
    CLASS CORE ;
    FOREIGN XOR3_0011 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.3600 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 3.2475 0.3075 3.3225 0.7350 ;
        RECT 3.0825 0.3075 3.2475 0.3825 ;
        RECT 3.0825 0.6600 3.2475 0.7350 ;
        RECT 3.0075 0.2175 3.0825 0.3825 ;
        RECT 3.0075 0.6600 3.0825 0.8325 ;
        END
    END Z
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 2.7750 0.1125 3.0900 0.1875 ;
        RECT 2.7000 0.1125 2.7750 0.4875 ;
        RECT 2.3850 0.4125 2.7000 0.4875 ;
        VIA 2.6850 0.4500 VIA12_square ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.2450 0.5625 1.7100 0.6375 ;
        VIA 1.3725 0.6000 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.1350 0.4125 0.6000 0.4875 ;
        VIA 0.3675 0.4500 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 3.3150 -0.0750 3.3600 0.0750 ;
        RECT 3.1950 -0.0750 3.3150 0.2325 ;
        RECT 2.8875 -0.0750 3.1950 0.0750 ;
        RECT 2.7825 -0.0750 2.8875 0.2550 ;
        RECT 1.8450 -0.0750 2.7825 0.0750 ;
        RECT 1.7250 -0.0750 1.8450 0.2400 ;
        RECT 1.4175 -0.0750 1.7250 0.0750 ;
        RECT 1.3050 -0.0750 1.4175 0.2550 ;
        RECT 0.3675 -0.0750 1.3050 0.0750 ;
        RECT 0.2625 -0.0750 0.3675 0.2550 ;
        RECT 0.0000 -0.0750 0.2625 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 3.3150 0.9750 3.3600 1.1250 ;
        RECT 3.1950 0.8100 3.3150 1.1250 ;
        RECT 2.8950 0.9750 3.1950 1.1250 ;
        RECT 2.7900 0.8100 2.8950 1.1250 ;
        RECT 1.8450 0.9750 2.7900 1.1250 ;
        RECT 1.7250 0.8175 1.8450 1.1250 ;
        RECT 1.4025 0.9750 1.7250 1.1250 ;
        RECT 1.3275 0.7875 1.4025 1.1250 ;
        RECT 0.3750 0.9750 1.3275 1.1250 ;
        RECT 0.2550 0.8250 0.3750 1.1250 ;
        RECT 0.0000 0.9750 0.2550 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 3.2250 0.1725 3.2850 0.2325 ;
        RECT 3.2250 0.8175 3.2850 0.8775 ;
        RECT 3.1125 0.4875 3.1725 0.5475 ;
        RECT 3.0150 0.2700 3.0750 0.3300 ;
        RECT 3.0150 0.7200 3.0750 0.7800 ;
        RECT 2.9100 0.4875 2.9700 0.5475 ;
        RECT 2.8050 0.1650 2.8650 0.2250 ;
        RECT 2.8050 0.8400 2.8650 0.9000 ;
        RECT 2.7000 0.4650 2.7600 0.5250 ;
        RECT 2.5950 0.1800 2.6550 0.2400 ;
        RECT 2.5950 0.6600 2.6550 0.7200 ;
        RECT 2.4900 0.4500 2.5500 0.5100 ;
        RECT 2.3850 0.1800 2.4450 0.2400 ;
        RECT 2.3850 0.8325 2.4450 0.8925 ;
        RECT 2.2800 0.5025 2.3400 0.5625 ;
        RECT 2.1750 0.1800 2.2350 0.2400 ;
        RECT 2.1750 0.8325 2.2350 0.8925 ;
        RECT 2.0700 0.6600 2.1300 0.7200 ;
        RECT 1.8600 0.3600 1.9200 0.4200 ;
        RECT 1.8600 0.6000 1.9200 0.6600 ;
        RECT 1.7550 0.1500 1.8150 0.2100 ;
        RECT 1.7550 0.8475 1.8150 0.9075 ;
        RECT 1.6500 0.5250 1.7100 0.5850 ;
        RECT 1.5450 0.1800 1.6050 0.2400 ;
        RECT 1.5450 0.8175 1.6050 0.8775 ;
        RECT 1.3350 0.1650 1.3950 0.2250 ;
        RECT 1.3350 0.8175 1.3950 0.8775 ;
        RECT 1.2300 0.5100 1.2900 0.5700 ;
        RECT 1.1250 0.1800 1.1850 0.2400 ;
        RECT 1.1250 0.7200 1.1850 0.7800 ;
        RECT 1.0200 0.4950 1.0800 0.5550 ;
        RECT 0.9150 0.1800 0.9750 0.2400 ;
        RECT 0.9150 0.8325 0.9750 0.8925 ;
        RECT 0.8025 0.6375 0.8625 0.6975 ;
        RECT 0.7050 0.1650 0.7650 0.2250 ;
        RECT 0.7050 0.8325 0.7650 0.8925 ;
        RECT 0.6000 0.3450 0.6600 0.4050 ;
        RECT 0.3900 0.4200 0.4500 0.4800 ;
        RECT 0.3900 0.6600 0.4500 0.7200 ;
        RECT 0.2850 0.1725 0.3450 0.2325 ;
        RECT 0.2850 0.8475 0.3450 0.9075 ;
        RECT 0.1875 0.4725 0.2475 0.5325 ;
        RECT 0.0750 0.2175 0.1350 0.2775 ;
        RECT 0.0750 0.8175 0.1350 0.8775 ;
        LAYER M1 ;
        RECT 2.9325 0.4575 3.1725 0.5775 ;
        RECT 2.8425 0.4575 2.9325 0.6825 ;
        RECT 2.6325 0.3300 2.7675 0.5700 ;
        RECT 2.4825 0.1500 2.6925 0.2550 ;
        RECT 2.5650 0.6450 2.6850 0.7500 ;
        RECT 2.0400 0.6450 2.5650 0.7350 ;
        RECT 2.4825 0.3450 2.5575 0.5400 ;
        RECT 2.3100 0.1500 2.4825 0.2700 ;
        RECT 1.6275 0.3450 2.4825 0.4200 ;
        RECT 2.0625 0.8100 2.4750 0.9000 ;
        RECT 1.9350 0.4950 2.3775 0.5700 ;
        RECT 1.9500 0.1500 2.2350 0.2700 ;
        RECT 1.8300 0.4950 1.9350 0.6900 ;
        RECT 1.6425 0.4950 1.8300 0.6150 ;
        RECT 1.5675 0.7950 1.6350 0.9000 ;
        RECT 1.5675 0.1500 1.6275 0.4200 ;
        RECT 1.5225 0.1500 1.5675 0.9000 ;
        RECT 1.4850 0.3450 1.5225 0.9000 ;
        RECT 1.3050 0.3675 1.4100 0.6825 ;
        RECT 1.1925 0.4875 1.3050 0.5925 ;
        RECT 1.1025 0.1500 1.2150 0.4125 ;
        RECT 1.1100 0.6675 1.2150 0.9000 ;
        RECT 1.0050 0.4875 1.1100 0.5925 ;
        RECT 1.0050 0.6675 1.1100 0.7425 ;
        RECT 0.9975 0.3375 1.1025 0.4125 ;
        RECT 0.4500 0.4875 1.0050 0.5625 ;
        RECT 0.6150 0.8175 1.0050 0.9000 ;
        RECT 0.8925 0.1500 0.9975 0.4125 ;
        RECT 0.5700 0.3375 0.8925 0.4125 ;
        RECT 0.1575 0.6375 0.8925 0.7200 ;
        RECT 0.4650 0.1500 0.7950 0.2550 ;
        RECT 0.3300 0.3675 0.4500 0.5625 ;
        RECT 0.1875 0.4425 0.3300 0.5625 ;
        RECT 0.1125 0.2100 0.1800 0.3300 ;
        RECT 0.1125 0.6375 0.1575 0.9000 ;
        RECT 0.0375 0.2100 0.1125 0.9000 ;
        LAYER VIA1 ;
        RECT 2.8425 0.5625 2.9175 0.6375 ;
        RECT 2.4075 0.6450 2.4825 0.7200 ;
        RECT 2.3475 0.1725 2.4225 0.2475 ;
        RECT 2.2575 0.8100 2.3325 0.8850 ;
        RECT 1.9950 0.1725 2.0700 0.2475 ;
        RECT 1.8450 0.4950 1.9200 0.5700 ;
        RECT 1.0950 0.3375 1.1700 0.4125 ;
        RECT 1.0500 0.6675 1.1250 0.7425 ;
        RECT 0.7275 0.8175 0.8025 0.8925 ;
        RECT 0.5775 0.1650 0.6525 0.2400 ;
        LAYER M2 ;
        RECT 2.8425 0.5625 2.9925 0.6375 ;
        RECT 2.7675 0.5625 2.8425 0.8850 ;
        RECT 2.1150 0.8100 2.7675 0.8850 ;
        RECT 2.2650 0.6450 2.5275 0.7200 ;
        RECT 2.2650 0.1725 2.4675 0.2475 ;
        RECT 2.1900 0.1725 2.2650 0.7200 ;
        RECT 2.0400 0.1725 2.1150 0.8850 ;
        RECT 1.9200 0.1725 2.0400 0.2475 ;
        RECT 1.8300 0.4125 1.9350 0.6150 ;
        RECT 1.4400 0.4125 1.8300 0.4875 ;
        RECT 1.3650 0.1650 1.4400 0.4875 ;
        RECT 0.8475 0.1650 1.3650 0.2400 ;
        RECT 1.1250 0.3375 1.2150 0.4125 ;
        RECT 1.0500 0.3375 1.1250 0.8250 ;
        RECT 0.7725 0.1650 0.8475 0.8925 ;
        RECT 0.5325 0.1650 0.7725 0.2400 ;
        RECT 0.6825 0.8175 0.7725 0.8925 ;
    END
END XOR3_0011


MACRO XOR3_0111
    CLASS CORE ;
    FOREIGN XOR3_0111 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.2000 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 3.5175 0.2625 3.8325 0.7275 ;
        VIA 3.6750 0.3225 VIA12_slot ;
        VIA 3.6750 0.6675 VIA12_slot ;
        END
    END Z
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 3.3375 0.6825 3.4425 0.7875 ;
        RECT 2.9625 0.7125 3.3375 0.7875 ;
        VIA 3.2550 0.7500 VIA12_square ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.2150 0.5625 1.6800 0.6375 ;
        VIA 1.3350 0.6000 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.1350 0.4125 0.6000 0.4875 ;
        VIA 0.3675 0.4500 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 4.1475 -0.0750 4.2000 0.0750 ;
        RECT 4.0425 -0.0750 4.1475 0.3000 ;
        RECT 3.7350 -0.0750 4.0425 0.0750 ;
        RECT 3.6150 -0.0750 3.7350 0.1950 ;
        RECT 3.3150 -0.0750 3.6150 0.0750 ;
        RECT 3.2250 -0.0750 3.3150 0.2925 ;
        RECT 2.2650 -0.0750 3.2250 0.0750 ;
        RECT 2.1450 -0.0750 2.2650 0.1875 ;
        RECT 1.4175 -0.0750 2.1450 0.0750 ;
        RECT 1.3050 -0.0750 1.4175 0.2550 ;
        RECT 0.3675 -0.0750 1.3050 0.0750 ;
        RECT 0.2625 -0.0750 0.3675 0.2550 ;
        RECT 0.0000 -0.0750 0.2625 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 4.1550 0.9750 4.2000 1.1250 ;
        RECT 4.0350 0.7725 4.1550 1.1250 ;
        RECT 3.7350 0.9750 4.0350 1.1250 ;
        RECT 3.6150 0.8175 3.7350 1.1250 ;
        RECT 3.3150 0.9750 3.6150 1.1250 ;
        RECT 3.1950 0.8625 3.3150 1.1250 ;
        RECT 1.8375 0.9750 3.1950 1.1250 ;
        RECT 1.7325 0.7500 1.8375 1.1250 ;
        RECT 1.4175 0.9750 1.7325 1.1250 ;
        RECT 1.3125 0.7875 1.4175 1.1250 ;
        RECT 0.3750 0.9750 1.3125 1.1250 ;
        RECT 0.2550 0.8250 0.3750 1.1250 ;
        RECT 0.0000 0.9750 0.2550 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 4.0650 0.2175 4.1250 0.2775 ;
        RECT 4.0650 0.7800 4.1250 0.8400 ;
        RECT 3.9525 0.4650 4.0125 0.5250 ;
        RECT 3.8550 0.2250 3.9150 0.2850 ;
        RECT 3.8550 0.6525 3.9150 0.7125 ;
        RECT 3.7500 0.4650 3.8100 0.5250 ;
        RECT 3.6450 0.1275 3.7050 0.1875 ;
        RECT 3.6450 0.8325 3.7050 0.8925 ;
        RECT 3.5400 0.4650 3.6000 0.5250 ;
        RECT 3.4350 0.2250 3.4950 0.2850 ;
        RECT 3.4350 0.6525 3.4950 0.7125 ;
        RECT 3.3300 0.4650 3.3900 0.5250 ;
        RECT 3.2250 0.2025 3.2850 0.2625 ;
        RECT 3.2250 0.8700 3.2850 0.9300 ;
        RECT 3.1200 0.4800 3.1800 0.5400 ;
        RECT 3.0150 0.1800 3.0750 0.2400 ;
        RECT 3.0150 0.8100 3.0750 0.8700 ;
        RECT 2.9100 0.4800 2.9700 0.5400 ;
        RECT 2.8050 0.1725 2.8650 0.2325 ;
        RECT 2.8050 0.8250 2.8650 0.8850 ;
        RECT 2.6925 0.4950 2.7525 0.5550 ;
        RECT 2.5950 0.1875 2.6550 0.2475 ;
        RECT 2.5950 0.8175 2.6550 0.8775 ;
        RECT 2.4900 0.6450 2.5500 0.7050 ;
        RECT 2.3850 0.2400 2.4450 0.3000 ;
        RECT 2.3850 0.8175 2.4450 0.8775 ;
        RECT 2.2800 0.4950 2.3400 0.5550 ;
        RECT 2.1750 0.1200 2.2350 0.1800 ;
        RECT 2.0700 0.4950 2.1300 0.5550 ;
        RECT 1.9650 0.2475 2.0250 0.3075 ;
        RECT 1.9650 0.7575 2.0250 0.8175 ;
        RECT 1.8600 0.4800 1.9200 0.5400 ;
        RECT 1.7550 0.7725 1.8150 0.8325 ;
        RECT 1.6500 0.4800 1.7100 0.5400 ;
        RECT 1.5450 0.2550 1.6050 0.3150 ;
        RECT 1.5450 0.8175 1.6050 0.8775 ;
        RECT 1.4475 0.4800 1.5075 0.5400 ;
        RECT 1.3350 0.1650 1.3950 0.2250 ;
        RECT 1.3350 0.8175 1.3950 0.8775 ;
        RECT 1.2300 0.4950 1.2900 0.5550 ;
        RECT 1.1250 0.1800 1.1850 0.2400 ;
        RECT 1.1250 0.7200 1.1850 0.7800 ;
        RECT 1.0200 0.4950 1.0800 0.5550 ;
        RECT 0.9150 0.1800 0.9750 0.2400 ;
        RECT 0.9150 0.8325 0.9750 0.8925 ;
        RECT 0.8025 0.6375 0.8625 0.6975 ;
        RECT 0.7050 0.1650 0.7650 0.2250 ;
        RECT 0.7050 0.8325 0.7650 0.8925 ;
        RECT 0.6000 0.3450 0.6600 0.4050 ;
        RECT 0.3900 0.4200 0.4500 0.4800 ;
        RECT 0.3900 0.6600 0.4500 0.7200 ;
        RECT 0.2850 0.1725 0.3450 0.2325 ;
        RECT 0.2850 0.8475 0.3450 0.9075 ;
        RECT 0.1875 0.4725 0.2475 0.5325 ;
        RECT 0.0750 0.2175 0.1350 0.2775 ;
        RECT 0.0750 0.8175 0.1350 0.8775 ;
        LAYER M1 ;
        RECT 3.9900 0.4425 4.0950 0.6825 ;
        RECT 3.2925 0.4425 3.9900 0.5475 ;
        RECT 3.8325 0.1950 3.9150 0.3675 ;
        RECT 3.4350 0.6225 3.9150 0.7425 ;
        RECT 3.5175 0.2775 3.8325 0.3675 ;
        RECT 3.4125 0.1950 3.5175 0.3675 ;
        RECT 3.2175 0.6450 3.3375 0.7875 ;
        RECT 3.1725 0.4650 3.2175 0.7875 ;
        RECT 3.1425 0.4650 3.1725 0.7050 ;
        RECT 3.0450 0.1500 3.1500 0.3900 ;
        RECT 3.0900 0.4650 3.1425 0.5700 ;
        RECT 3.0675 0.7800 3.0975 0.9000 ;
        RECT 2.9925 0.6450 3.0675 0.9000 ;
        RECT 2.7825 0.1500 3.0450 0.2550 ;
        RECT 2.9700 0.4650 3.0150 0.5700 ;
        RECT 2.4600 0.6450 2.9925 0.7200 ;
        RECT 2.8875 0.3300 2.9700 0.5700 ;
        RECT 2.5425 0.7950 2.9175 0.9000 ;
        RECT 2.7825 0.3300 2.8875 0.4050 ;
        RECT 2.5875 0.4800 2.7825 0.5700 ;
        RECT 2.6550 0.1500 2.6775 0.2850 ;
        RECT 2.5275 0.1500 2.6550 0.3900 ;
        RECT 2.4300 0.4650 2.5875 0.5700 ;
        RECT 2.3475 0.7950 2.4675 0.9000 ;
        RECT 2.3775 0.1950 2.4525 0.3375 ;
        RECT 2.0400 0.2625 2.3775 0.3375 ;
        RECT 2.1300 0.4125 2.3550 0.5850 ;
        RECT 2.2050 0.6600 2.3475 0.9000 ;
        RECT 2.0550 0.4125 2.1300 0.8400 ;
        RECT 1.9425 0.7350 2.0550 0.8400 ;
        RECT 1.9500 0.2175 2.0400 0.3375 ;
        RECT 1.4475 0.4500 1.9500 0.5700 ;
        RECT 1.5150 0.1650 1.7625 0.3750 ;
        RECT 1.4925 0.6600 1.6575 0.9000 ;
        RECT 1.2900 0.3600 1.3725 0.6825 ;
        RECT 1.1925 0.4875 1.2900 0.5925 ;
        RECT 1.1025 0.1500 1.2150 0.4125 ;
        RECT 1.1100 0.6675 1.2150 0.9000 ;
        RECT 1.0050 0.4875 1.1100 0.5925 ;
        RECT 1.0050 0.6675 1.1100 0.7425 ;
        RECT 0.9975 0.3375 1.1025 0.4125 ;
        RECT 0.4500 0.4875 1.0050 0.5625 ;
        RECT 0.6150 0.8175 1.0050 0.9000 ;
        RECT 0.8925 0.1500 0.9975 0.4125 ;
        RECT 0.5700 0.3375 0.8925 0.4125 ;
        RECT 0.1575 0.6375 0.8925 0.7200 ;
        RECT 0.4650 0.1500 0.7950 0.2550 ;
        RECT 0.3300 0.3675 0.4500 0.5625 ;
        RECT 0.1875 0.4425 0.3300 0.5625 ;
        RECT 0.1125 0.2100 0.1800 0.3300 ;
        RECT 0.1125 0.6375 0.1575 0.9000 ;
        RECT 0.0375 0.2100 0.1125 0.9000 ;
        LAYER VIA1 ;
        RECT 3.9900 0.5625 4.0650 0.6375 ;
        RECT 3.3300 0.4575 3.4050 0.5325 ;
        RECT 3.0600 0.2775 3.1350 0.3525 ;
        RECT 2.8275 0.3300 2.9025 0.4050 ;
        RECT 2.7525 0.6450 2.8275 0.7200 ;
        RECT 2.5800 0.8100 2.6550 0.8850 ;
        RECT 2.5650 0.1650 2.6400 0.2400 ;
        RECT 2.4675 0.4800 2.5425 0.5550 ;
        RECT 2.2350 0.7125 2.3100 0.7875 ;
        RECT 2.1225 0.4125 2.1975 0.4875 ;
        RECT 1.8000 0.4650 1.8750 0.5400 ;
        RECT 1.6350 0.2625 1.7100 0.3375 ;
        RECT 1.5375 0.7125 1.6125 0.7875 ;
        RECT 1.1250 0.7125 1.2000 0.7875 ;
        RECT 1.0950 0.3375 1.1700 0.4125 ;
        RECT 0.7275 0.8175 0.8025 0.8925 ;
        RECT 0.5775 0.1650 0.6525 0.2400 ;
        LAYER M2 ;
        RECT 3.9975 0.5625 4.1400 0.6375 ;
        RECT 3.9225 0.5625 3.9975 0.9375 ;
        RECT 2.6550 0.8625 3.9225 0.9375 ;
        RECT 3.3225 0.4200 3.4200 0.5700 ;
        RECT 3.2475 0.1125 3.3225 0.5700 ;
        RECT 2.7000 0.1125 3.2475 0.1875 ;
        RECT 3.0675 0.2625 3.1725 0.3675 ;
        RECT 2.9925 0.2625 3.0675 0.6375 ;
        RECT 2.8425 0.5625 2.9925 0.6375 ;
        RECT 2.8125 0.2925 2.9175 0.4425 ;
        RECT 2.7375 0.5625 2.8425 0.7650 ;
        RECT 2.2725 0.3150 2.8125 0.3900 ;
        RECT 2.6250 0.1125 2.7000 0.2400 ;
        RECT 2.5800 0.7650 2.6550 0.9375 ;
        RECT 2.4900 0.1650 2.6250 0.2400 ;
        RECT 2.4375 0.4650 2.5800 0.5700 ;
        RECT 2.3475 0.4650 2.4375 0.6375 ;
        RECT 1.4625 0.7125 2.3850 0.7875 ;
        RECT 1.8750 0.5625 2.3475 0.6375 ;
        RECT 2.1975 0.3150 2.2725 0.4875 ;
        RECT 2.0250 0.4125 2.1975 0.4875 ;
        RECT 1.9500 0.2625 2.0250 0.4875 ;
        RECT 1.5600 0.2625 1.9500 0.3375 ;
        RECT 1.8000 0.4125 1.8750 0.6375 ;
        RECT 1.4400 0.4125 1.8000 0.4875 ;
        RECT 1.3650 0.1650 1.4400 0.4875 ;
        RECT 0.8475 0.1650 1.3650 0.2400 ;
        RECT 1.0950 0.7125 1.2750 0.7875 ;
        RECT 1.0950 0.3375 1.2150 0.4125 ;
        RECT 1.0200 0.3375 1.0950 0.7875 ;
        RECT 0.7725 0.1650 0.8475 0.8925 ;
        RECT 0.5325 0.1650 0.7725 0.2400 ;
        RECT 0.6825 0.8175 0.7725 0.8925 ;
    END
END XOR3_0111


MACRO XOR3_1000
    CLASS CORE ;
    FOREIGN XOR3_1000 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.7700 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 7.0875 0.3075 7.4025 0.7425 ;
        VIA 7.2450 0.3750 VIA12_slot ;
        VIA 7.2450 0.6750 VIA12_slot ;
        END
    END Z
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 5.5425 0.4125 6.0975 0.4875 ;
        RECT 5.4375 0.4125 5.5425 0.6075 ;
        VIA 5.9775 0.4500 VIA12_square ;
        VIA 5.4900 0.5175 VIA12_square ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.9000 0.4350 1.0125 0.6375 ;
        RECT 0.3900 0.5625 0.9000 0.6375 ;
        VIA 0.9600 0.5175 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 2.1825 0.4125 2.7375 0.4875 ;
        RECT 2.0775 0.4125 2.1825 0.6075 ;
        VIA 2.6175 0.4500 VIA12_square ;
        VIA 2.1300 0.5175 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 5.8500 -0.0750 7.7700 0.0750 ;
        RECT 5.7000 -0.0750 5.8500 0.2175 ;
        RECT 5.4150 -0.0750 5.7000 0.0750 ;
        RECT 5.2950 -0.0750 5.4150 0.2250 ;
        RECT 4.9950 -0.0750 5.2950 0.0750 ;
        RECT 4.8750 -0.0750 4.9950 0.2325 ;
        RECT 4.5750 -0.0750 4.8750 0.0750 ;
        RECT 4.4550 -0.0750 4.5750 0.2325 ;
        RECT 2.4900 -0.0750 4.4550 0.0750 ;
        RECT 2.3400 -0.0750 2.4900 0.2175 ;
        RECT 2.0550 -0.0750 2.3400 0.0750 ;
        RECT 1.9350 -0.0750 2.0550 0.2250 ;
        RECT 1.6350 -0.0750 1.9350 0.0750 ;
        RECT 1.5150 -0.0750 1.6350 0.2325 ;
        RECT 1.2150 -0.0750 1.5150 0.0750 ;
        RECT 1.0950 -0.0750 1.2150 0.2325 ;
        RECT 0.7950 -0.0750 1.0950 0.0750 ;
        RECT 0.6750 -0.0750 0.7950 0.2325 ;
        RECT 0.3675 -0.0750 0.6750 0.0750 ;
        RECT 0.2625 -0.0750 0.3675 0.2325 ;
        RECT 0.0000 -0.0750 0.2625 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 5.8350 0.9750 7.7700 1.1250 ;
        RECT 5.7150 0.8325 5.8350 1.1250 ;
        RECT 5.4300 0.9750 5.7150 1.1250 ;
        RECT 5.2800 0.8325 5.4300 1.1250 ;
        RECT 4.9950 0.9750 5.2800 1.1250 ;
        RECT 4.8750 0.8400 4.9950 1.1250 ;
        RECT 4.5750 0.9750 4.8750 1.1250 ;
        RECT 4.4550 0.8250 4.5750 1.1250 ;
        RECT 2.4750 0.9750 4.4550 1.1250 ;
        RECT 2.3550 0.8325 2.4750 1.1250 ;
        RECT 2.0700 0.9750 2.3550 1.1250 ;
        RECT 1.9200 0.8325 2.0700 1.1250 ;
        RECT 1.6350 0.9750 1.9200 1.1250 ;
        RECT 1.5150 0.8400 1.6350 1.1250 ;
        RECT 1.2150 0.9750 1.5150 1.1250 ;
        RECT 1.0950 0.8400 1.2150 1.1250 ;
        RECT 0.7950 0.9750 1.0950 1.1250 ;
        RECT 0.6750 0.8400 0.7950 1.1250 ;
        RECT 0.3750 0.9750 0.6750 1.1250 ;
        RECT 0.2550 0.8400 0.3750 1.1250 ;
        RECT 0.0000 0.9750 0.2550 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 7.6350 0.3075 7.6950 0.3675 ;
        RECT 7.6350 0.6750 7.6950 0.7350 ;
        RECT 7.5300 0.4950 7.5900 0.5550 ;
        RECT 7.4250 0.1575 7.4850 0.2175 ;
        RECT 7.4250 0.8325 7.4850 0.8925 ;
        RECT 7.3200 0.4950 7.3800 0.5550 ;
        RECT 7.2150 0.3225 7.2750 0.3825 ;
        RECT 7.2150 0.6750 7.2750 0.7350 ;
        RECT 7.1100 0.4950 7.1700 0.5550 ;
        RECT 7.0050 0.1575 7.0650 0.2175 ;
        RECT 7.0050 0.8325 7.0650 0.8925 ;
        RECT 6.9000 0.4950 6.9600 0.5550 ;
        RECT 6.7950 0.2625 6.8550 0.3225 ;
        RECT 6.7950 0.6750 6.8550 0.7350 ;
        RECT 6.6900 0.4800 6.7500 0.5400 ;
        RECT 6.5850 0.3000 6.6450 0.3600 ;
        RECT 6.5850 0.6675 6.6450 0.7275 ;
        RECT 6.4800 0.4800 6.5400 0.5400 ;
        RECT 6.3750 0.1575 6.4350 0.2175 ;
        RECT 6.3750 0.8325 6.4350 0.8925 ;
        RECT 6.2700 0.4800 6.3300 0.5400 ;
        RECT 6.1650 0.3000 6.2250 0.3600 ;
        RECT 6.1650 0.6825 6.2250 0.7425 ;
        RECT 6.0600 0.4800 6.1200 0.5400 ;
        RECT 5.9550 0.1875 6.0150 0.2475 ;
        RECT 5.9550 0.8025 6.0150 0.8625 ;
        RECT 5.7450 0.1575 5.8050 0.2175 ;
        RECT 5.7450 0.8325 5.8050 0.8925 ;
        RECT 5.6400 0.4875 5.7000 0.5475 ;
        RECT 5.5350 0.3075 5.5950 0.3675 ;
        RECT 5.5350 0.6900 5.5950 0.7500 ;
        RECT 5.4300 0.4875 5.4900 0.5475 ;
        RECT 5.3250 0.1425 5.3850 0.2025 ;
        RECT 5.3250 0.8325 5.3850 0.8925 ;
        RECT 5.2200 0.4875 5.2800 0.5475 ;
        RECT 5.1150 0.2925 5.1750 0.3525 ;
        RECT 5.1150 0.7200 5.1750 0.7800 ;
        RECT 5.0100 0.4875 5.0700 0.5475 ;
        RECT 4.9050 0.1650 4.9650 0.2250 ;
        RECT 4.9050 0.8475 4.9650 0.9075 ;
        RECT 4.8000 0.4875 4.8600 0.5475 ;
        RECT 4.6950 0.2925 4.7550 0.3525 ;
        RECT 4.6950 0.7350 4.7550 0.7950 ;
        RECT 4.5900 0.4875 4.6500 0.5475 ;
        RECT 4.4850 0.1650 4.5450 0.2250 ;
        RECT 4.4850 0.8325 4.5450 0.8925 ;
        RECT 4.2750 0.3075 4.3350 0.3675 ;
        RECT 4.2750 0.6750 4.3350 0.7350 ;
        RECT 4.1700 0.4950 4.2300 0.5550 ;
        RECT 4.0650 0.1575 4.1250 0.2175 ;
        RECT 4.0650 0.8325 4.1250 0.8925 ;
        RECT 3.9600 0.4950 4.0200 0.5550 ;
        RECT 3.8550 0.3225 3.9150 0.3825 ;
        RECT 3.8550 0.6750 3.9150 0.7350 ;
        RECT 3.7500 0.4950 3.8100 0.5550 ;
        RECT 3.6450 0.1575 3.7050 0.2175 ;
        RECT 3.6450 0.8325 3.7050 0.8925 ;
        RECT 3.5400 0.4950 3.6000 0.5550 ;
        RECT 3.4350 0.2625 3.4950 0.3225 ;
        RECT 3.4350 0.6750 3.4950 0.7350 ;
        RECT 3.3300 0.4800 3.3900 0.5400 ;
        RECT 3.2250 0.3000 3.2850 0.3600 ;
        RECT 3.2250 0.6675 3.2850 0.7275 ;
        RECT 3.1200 0.4800 3.1800 0.5400 ;
        RECT 3.0150 0.1575 3.0750 0.2175 ;
        RECT 3.0150 0.8325 3.0750 0.8925 ;
        RECT 2.9100 0.4800 2.9700 0.5400 ;
        RECT 2.8050 0.3000 2.8650 0.3600 ;
        RECT 2.8050 0.6825 2.8650 0.7425 ;
        RECT 2.7000 0.4800 2.7600 0.5400 ;
        RECT 2.5950 0.1875 2.6550 0.2475 ;
        RECT 2.5950 0.8025 2.6550 0.8625 ;
        RECT 2.3850 0.1575 2.4450 0.2175 ;
        RECT 2.3850 0.8325 2.4450 0.8925 ;
        RECT 2.2800 0.4875 2.3400 0.5475 ;
        RECT 2.1750 0.3075 2.2350 0.3675 ;
        RECT 2.1750 0.6900 2.2350 0.7500 ;
        RECT 2.0700 0.4875 2.1300 0.5475 ;
        RECT 1.9650 0.1425 2.0250 0.2025 ;
        RECT 1.9650 0.8325 2.0250 0.8925 ;
        RECT 1.8600 0.4875 1.9200 0.5475 ;
        RECT 1.7550 0.2925 1.8150 0.3525 ;
        RECT 1.7550 0.7200 1.8150 0.7800 ;
        RECT 1.6500 0.4875 1.7100 0.5475 ;
        RECT 1.5450 0.1650 1.6050 0.2250 ;
        RECT 1.5450 0.8475 1.6050 0.9075 ;
        RECT 1.4400 0.4875 1.5000 0.5475 ;
        RECT 1.3350 0.2925 1.3950 0.3525 ;
        RECT 1.3350 0.7350 1.3950 0.7950 ;
        RECT 1.2300 0.4875 1.2900 0.5475 ;
        RECT 1.1250 0.1650 1.1850 0.2250 ;
        RECT 1.1250 0.8475 1.1850 0.9075 ;
        RECT 1.0200 0.4875 1.0800 0.5475 ;
        RECT 0.9150 0.2925 0.9750 0.3525 ;
        RECT 0.9150 0.7350 0.9750 0.7950 ;
        RECT 0.8100 0.4875 0.8700 0.5475 ;
        RECT 0.7050 0.1650 0.7650 0.2250 ;
        RECT 0.7050 0.8475 0.7650 0.9075 ;
        RECT 0.6000 0.4875 0.6600 0.5475 ;
        RECT 0.4950 0.2925 0.5550 0.3525 ;
        RECT 0.4950 0.7350 0.5550 0.7950 ;
        RECT 0.3900 0.4875 0.4500 0.5475 ;
        RECT 0.2850 0.1500 0.3450 0.2100 ;
        RECT 0.2850 0.8475 0.3450 0.9075 ;
        RECT 0.1800 0.4875 0.2400 0.5475 ;
        RECT 0.0750 0.2925 0.1350 0.3525 ;
        RECT 0.0750 0.7350 0.1350 0.7950 ;
        LAYER M1 ;
        RECT 7.6050 0.2775 7.7250 0.4125 ;
        RECT 7.6200 0.6375 7.7025 0.7875 ;
        RECT 7.0200 0.4875 7.6500 0.5625 ;
        RECT 7.0875 0.6375 7.6200 0.7350 ;
        RECT 7.0875 0.3075 7.6050 0.4125 ;
        RECT 7.1325 0.1500 7.5375 0.2250 ;
        RECT 7.0875 0.8250 7.5150 0.9000 ;
        RECT 6.9675 0.1500 7.1325 0.2325 ;
        RECT 6.8625 0.3075 7.0875 0.3825 ;
        RECT 6.8175 0.6600 7.0875 0.7350 ;
        RECT 6.9225 0.8175 7.0875 0.9000 ;
        RECT 6.8250 0.4575 7.0200 0.5850 ;
        RECT 6.7875 0.1500 6.8625 0.3825 ;
        RECT 6.7425 0.6600 6.8175 0.9000 ;
        RECT 6.0300 0.1500 6.7875 0.2250 ;
        RECT 6.6450 0.4500 6.7500 0.5700 ;
        RECT 6.0225 0.8250 6.7425 0.9000 ;
        RECT 6.1350 0.3000 6.6750 0.3750 ;
        RECT 6.5025 0.6450 6.6675 0.7500 ;
        RECT 6.0300 0.4500 6.6450 0.5400 ;
        RECT 6.1350 0.6750 6.5025 0.7500 ;
        RECT 5.9250 0.1500 6.0300 0.2850 ;
        RECT 5.9250 0.3750 6.0300 0.5400 ;
        RECT 5.9475 0.7575 6.0225 0.9000 ;
        RECT 5.7750 0.3075 5.8500 0.7575 ;
        RECT 5.4975 0.3075 5.7750 0.3825 ;
        RECT 5.4300 0.6525 5.7750 0.7575 ;
        RECT 5.3925 0.4575 5.7000 0.5775 ;
        RECT 4.5300 0.4725 5.3100 0.5775 ;
        RECT 5.1825 0.3075 5.2725 0.3825 ;
        RECT 5.1075 0.2625 5.1825 0.3825 ;
        RECT 5.1075 0.6825 5.1825 0.8175 ;
        RECT 4.7625 0.3075 5.1075 0.3825 ;
        RECT 4.7625 0.6825 5.1075 0.7575 ;
        RECT 4.6875 0.2250 4.7625 0.3825 ;
        RECT 4.6875 0.6825 4.7625 0.8400 ;
        RECT 4.4550 0.3075 4.5300 0.7350 ;
        RECT 3.5025 0.3075 4.4550 0.3825 ;
        RECT 3.4575 0.6600 4.4550 0.7350 ;
        RECT 3.6600 0.4875 4.2900 0.5625 ;
        RECT 3.7725 0.1500 4.1775 0.2250 ;
        RECT 3.7275 0.8250 4.1550 0.9000 ;
        RECT 3.6075 0.1500 3.7725 0.2325 ;
        RECT 3.5625 0.8175 3.7275 0.9000 ;
        RECT 3.4650 0.4575 3.6600 0.5850 ;
        RECT 3.4275 0.1500 3.5025 0.3825 ;
        RECT 3.3825 0.6600 3.4575 0.9000 ;
        RECT 2.6700 0.1500 3.4275 0.2250 ;
        RECT 3.2850 0.4500 3.3900 0.5700 ;
        RECT 2.6625 0.8250 3.3825 0.9000 ;
        RECT 2.7750 0.3000 3.3150 0.3750 ;
        RECT 3.1425 0.6450 3.3075 0.7500 ;
        RECT 2.6700 0.4500 3.2850 0.5400 ;
        RECT 2.7750 0.6750 3.1425 0.7500 ;
        RECT 2.5650 0.1500 2.6700 0.2850 ;
        RECT 2.5650 0.3750 2.6700 0.5400 ;
        RECT 2.5875 0.7575 2.6625 0.9000 ;
        RECT 2.4150 0.3075 2.4900 0.7575 ;
        RECT 2.1375 0.3075 2.4150 0.3825 ;
        RECT 2.0700 0.6525 2.4150 0.7575 ;
        RECT 2.0325 0.4575 2.3400 0.5775 ;
        RECT 1.7925 0.4725 1.9500 0.5775 ;
        RECT 1.8225 0.3075 1.9125 0.3825 ;
        RECT 1.8225 0.6600 1.9125 0.7350 ;
        RECT 1.7475 0.2625 1.8225 0.3825 ;
        RECT 1.7475 0.6600 1.8225 0.8175 ;
        RECT 1.2300 0.4575 1.7925 0.5775 ;
        RECT 1.4025 0.3075 1.7475 0.3825 ;
        RECT 1.4025 0.6600 1.7475 0.7350 ;
        RECT 1.3275 0.2250 1.4025 0.3825 ;
        RECT 1.3275 0.6600 1.4025 0.8400 ;
        RECT 1.1550 0.3075 1.2300 0.7575 ;
        RECT 0.9825 0.3075 1.1550 0.3825 ;
        RECT 0.9825 0.6825 1.1550 0.7575 ;
        RECT 0.1500 0.4575 1.0800 0.5775 ;
        RECT 0.9075 0.2325 0.9825 0.3825 ;
        RECT 0.9075 0.6825 0.9825 0.8400 ;
        RECT 0.5625 0.3075 0.9075 0.3825 ;
        RECT 0.5625 0.6825 0.9075 0.7575 ;
        RECT 0.4875 0.2325 0.5625 0.3825 ;
        RECT 0.4875 0.6825 0.5625 0.8400 ;
        RECT 0.1425 0.3075 0.4875 0.3825 ;
        RECT 0.1425 0.6825 0.4875 0.7575 ;
        RECT 0.0675 0.2325 0.1425 0.3825 ;
        RECT 0.0675 0.6825 0.1425 0.8400 ;
        LAYER VIA1 ;
        RECT 7.0125 0.1575 7.0875 0.2325 ;
        RECT 6.9675 0.8175 7.0425 0.8925 ;
        RECT 6.8625 0.4800 6.9375 0.5550 ;
        RECT 6.5475 0.6675 6.6225 0.7425 ;
        RECT 6.3225 0.3000 6.3975 0.3750 ;
        RECT 5.7750 0.5625 5.8500 0.6375 ;
        RECT 5.1450 0.3075 5.2200 0.3825 ;
        RECT 4.9425 0.4875 5.0175 0.5625 ;
        RECT 4.7775 0.3075 4.8525 0.3825 ;
        RECT 4.7775 0.6825 4.8525 0.7575 ;
        RECT 3.6525 0.1575 3.7275 0.2325 ;
        RECT 3.6075 0.8175 3.6825 0.8925 ;
        RECT 3.5025 0.4725 3.5775 0.5475 ;
        RECT 3.1875 0.6675 3.2625 0.7425 ;
        RECT 3.1650 0.3000 3.2400 0.3750 ;
        RECT 2.4150 0.5625 2.4900 0.6375 ;
        RECT 1.7475 0.3075 1.8225 0.3825 ;
        RECT 1.7475 0.6600 1.8225 0.7350 ;
        RECT 1.5375 0.4800 1.6125 0.5550 ;
        LAYER M2 ;
        RECT 6.9675 0.1125 7.1325 0.2325 ;
        RECT 6.9225 0.8175 7.0875 0.9375 ;
        RECT 5.0175 0.1125 6.9675 0.1875 ;
        RECT 6.8625 0.4275 6.9375 0.6225 ;
        RECT 4.8675 0.8625 6.9225 0.9375 ;
        RECT 6.6375 0.4275 6.8625 0.5025 ;
        RECT 6.5325 0.6225 6.6450 0.7875 ;
        RECT 6.5625 0.4275 6.6375 0.5475 ;
        RECT 6.4575 0.4725 6.5625 0.5475 ;
        RECT 5.0175 0.7125 6.5325 0.7875 ;
        RECT 6.3825 0.4725 6.4575 0.6375 ;
        RECT 6.2775 0.2625 6.4425 0.3900 ;
        RECT 5.7150 0.5625 6.3825 0.6375 ;
        RECT 5.2350 0.2625 6.2775 0.3375 ;
        RECT 5.1300 0.2625 5.2350 0.4275 ;
        RECT 4.9425 0.1125 5.0175 0.7875 ;
        RECT 4.7625 0.2625 4.8675 0.9375 ;
        RECT 3.8100 0.3150 3.8850 0.8925 ;
        RECT 3.3525 0.3150 3.8100 0.3900 ;
        RECT 3.6375 0.8175 3.8100 0.8925 ;
        RECT 3.5550 0.1575 3.7725 0.2325 ;
        RECT 3.5625 0.8175 3.6375 0.9375 ;
        RECT 3.0975 0.4725 3.6300 0.5475 ;
        RECT 1.6125 0.8625 3.5625 0.9375 ;
        RECT 3.4800 0.1125 3.5550 0.2325 ;
        RECT 1.8225 0.1125 3.4800 0.1875 ;
        RECT 3.3000 0.3000 3.3525 0.3900 ;
        RECT 3.1050 0.3000 3.3000 0.3750 ;
        RECT 3.1725 0.6225 3.2850 0.7875 ;
        RECT 1.8225 0.7125 3.1725 0.7875 ;
        RECT 3.0225 0.4725 3.0975 0.6375 ;
        RECT 2.3550 0.5625 3.0225 0.6375 ;
        RECT 1.7475 0.1125 1.8225 0.7875 ;
        RECT 1.5375 0.3075 1.6125 0.9375 ;
        RECT 1.3875 0.3075 1.5375 0.3825 ;
    END
END XOR3_1000


MACRO XOR3_1010
    CLASS CORE ;
    FOREIGN XOR3_1010 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.1500 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 3.0375 0.2175 3.1125 0.8325 ;
        RECT 3.0075 0.2175 3.0375 0.3825 ;
        RECT 3.0075 0.6675 3.0375 0.8325 ;
        END
    END Z
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 2.3250 0.4125 2.7900 0.4875 ;
        VIA 2.7000 0.4500 VIA12_square ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.2450 0.5625 1.7100 0.6375 ;
        VIA 1.3725 0.6000 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.1350 0.4125 0.6000 0.4875 ;
        VIA 0.3675 0.4500 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 2.8800 -0.0750 3.1500 0.0750 ;
        RECT 2.7750 -0.0750 2.8800 0.2100 ;
        RECT 1.8450 -0.0750 2.7750 0.0750 ;
        RECT 1.7250 -0.0750 1.8450 0.2400 ;
        RECT 1.4175 -0.0750 1.7250 0.0750 ;
        RECT 1.3050 -0.0750 1.4175 0.2550 ;
        RECT 0.3675 -0.0750 1.3050 0.0750 ;
        RECT 0.2625 -0.0750 0.3675 0.2550 ;
        RECT 0.0000 -0.0750 0.2625 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 2.8950 0.9750 3.1500 1.1250 ;
        RECT 2.7750 0.8700 2.8950 1.1250 ;
        RECT 1.8450 0.9750 2.7750 1.1250 ;
        RECT 1.7250 0.8175 1.8450 1.1250 ;
        RECT 1.4025 0.9750 1.7250 1.1250 ;
        RECT 1.3275 0.7875 1.4025 1.1250 ;
        RECT 0.3750 0.9750 1.3275 1.1250 ;
        RECT 0.2550 0.8250 0.3750 1.1250 ;
        RECT 0.0000 0.9750 0.2550 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 3.0150 0.2700 3.0750 0.3300 ;
        RECT 3.0150 0.7200 3.0750 0.7800 ;
        RECT 2.9025 0.4950 2.9625 0.5550 ;
        RECT 2.8050 0.1200 2.8650 0.1800 ;
        RECT 2.8050 0.8700 2.8650 0.9300 ;
        RECT 2.7000 0.4650 2.7600 0.5250 ;
        RECT 2.5950 0.1800 2.6550 0.2400 ;
        RECT 2.5950 0.7050 2.6550 0.7650 ;
        RECT 2.4825 0.4500 2.5425 0.5100 ;
        RECT 2.3850 0.1800 2.4450 0.2400 ;
        RECT 2.3850 0.8325 2.4450 0.8925 ;
        RECT 2.2725 0.5025 2.3325 0.5625 ;
        RECT 2.1750 0.1800 2.2350 0.2400 ;
        RECT 2.1750 0.8325 2.2350 0.8925 ;
        RECT 2.0700 0.6600 2.1300 0.7200 ;
        RECT 1.8600 0.3600 1.9200 0.4200 ;
        RECT 1.8600 0.6300 1.9200 0.6900 ;
        RECT 1.7550 0.1500 1.8150 0.2100 ;
        RECT 1.7550 0.8475 1.8150 0.9075 ;
        RECT 1.6500 0.5250 1.7100 0.5850 ;
        RECT 1.5450 0.1800 1.6050 0.2400 ;
        RECT 1.5450 0.8175 1.6050 0.8775 ;
        RECT 1.3350 0.1650 1.3950 0.2250 ;
        RECT 1.3350 0.8175 1.3950 0.8775 ;
        RECT 1.2300 0.5100 1.2900 0.5700 ;
        RECT 1.1250 0.1800 1.1850 0.2400 ;
        RECT 1.1250 0.7200 1.1850 0.7800 ;
        RECT 1.0200 0.4950 1.0800 0.5550 ;
        RECT 0.9150 0.1800 0.9750 0.2400 ;
        RECT 0.9150 0.8325 0.9750 0.8925 ;
        RECT 0.8025 0.6375 0.8625 0.6975 ;
        RECT 0.7050 0.1650 0.7650 0.2250 ;
        RECT 0.7050 0.8325 0.7650 0.8925 ;
        RECT 0.6000 0.3450 0.6600 0.4050 ;
        RECT 0.3900 0.4200 0.4500 0.4800 ;
        RECT 0.3900 0.6600 0.4500 0.7200 ;
        RECT 0.2850 0.1725 0.3450 0.2325 ;
        RECT 0.2850 0.8475 0.3450 0.9075 ;
        RECT 0.1875 0.4725 0.2475 0.5325 ;
        RECT 0.0750 0.2175 0.1350 0.2775 ;
        RECT 0.0750 0.8175 0.1350 0.8775 ;
        LAYER M1 ;
        RECT 2.9175 0.4650 2.9625 0.6075 ;
        RECT 2.8425 0.4650 2.9175 0.7950 ;
        RECT 2.7300 0.6300 2.8425 0.7950 ;
        RECT 2.6250 0.3300 2.7675 0.5550 ;
        RECT 2.4825 0.1500 2.6925 0.2550 ;
        RECT 2.5800 0.6450 2.6550 0.8325 ;
        RECT 2.0400 0.6450 2.5800 0.7350 ;
        RECT 2.4750 0.3450 2.5500 0.5400 ;
        RECT 2.3775 0.1500 2.4825 0.2700 ;
        RECT 1.6275 0.3450 2.4750 0.4200 ;
        RECT 2.0625 0.8100 2.4750 0.9000 ;
        RECT 1.9350 0.4950 2.3700 0.5700 ;
        RECT 1.9200 0.1500 2.3025 0.2700 ;
        RECT 1.8300 0.4950 1.9350 0.7200 ;
        RECT 1.6425 0.4950 1.8300 0.6150 ;
        RECT 1.5675 0.7950 1.6350 0.9000 ;
        RECT 1.5675 0.1500 1.6275 0.4200 ;
        RECT 1.5225 0.1500 1.5675 0.9000 ;
        RECT 1.4850 0.3450 1.5225 0.9000 ;
        RECT 1.3050 0.3675 1.4100 0.6825 ;
        RECT 1.1925 0.4875 1.3050 0.5925 ;
        RECT 1.1025 0.1500 1.2150 0.4125 ;
        RECT 1.1100 0.6675 1.2150 0.9000 ;
        RECT 1.0050 0.4875 1.1100 0.5925 ;
        RECT 1.0050 0.6675 1.1100 0.7425 ;
        RECT 0.9975 0.3375 1.1025 0.4125 ;
        RECT 0.4500 0.4875 1.0050 0.5625 ;
        RECT 0.6150 0.8175 1.0050 0.9000 ;
        RECT 0.8925 0.1500 0.9975 0.4125 ;
        RECT 0.5700 0.3375 0.8925 0.4125 ;
        RECT 0.1575 0.6375 0.8925 0.7200 ;
        RECT 0.4650 0.1500 0.7950 0.2550 ;
        RECT 0.3300 0.3675 0.4500 0.5625 ;
        RECT 0.1875 0.4425 0.3300 0.5625 ;
        RECT 0.1125 0.2100 0.1800 0.3300 ;
        RECT 0.1125 0.6375 0.1575 0.9000 ;
        RECT 0.0375 0.2100 0.1125 0.9000 ;
        LAYER VIA1 ;
        RECT 2.7750 0.7125 2.8500 0.7875 ;
        RECT 2.5275 0.1725 2.6025 0.2475 ;
        RECT 2.3775 0.6450 2.4525 0.7200 ;
        RECT 2.1075 0.8100 2.1825 0.8850 ;
        RECT 1.9650 0.1725 2.0400 0.2475 ;
        RECT 1.8300 0.4950 1.9050 0.5700 ;
        RECT 1.0950 0.3375 1.1700 0.4125 ;
        RECT 1.0500 0.6675 1.1250 0.7425 ;
        RECT 0.7275 0.8175 0.8025 0.8925 ;
        RECT 0.5775 0.1650 0.6525 0.2400 ;
        LAYER M2 ;
        RECT 2.7225 0.7125 2.9025 0.7875 ;
        RECT 2.6475 0.7125 2.7225 0.8850 ;
        RECT 2.2050 0.1725 2.6550 0.2475 ;
        RECT 2.0550 0.8100 2.6475 0.8850 ;
        RECT 2.2050 0.6450 2.4975 0.7200 ;
        RECT 2.1300 0.1725 2.2050 0.7200 ;
        RECT 1.9800 0.1350 2.0550 0.8850 ;
        RECT 1.9500 0.1350 1.9800 0.2850 ;
        RECT 1.8300 0.3675 1.9050 0.6525 ;
        RECT 1.8000 0.3675 1.8300 0.4425 ;
        RECT 1.7250 0.1650 1.8000 0.4425 ;
        RECT 0.8475 0.1650 1.7250 0.2400 ;
        RECT 1.1250 0.3375 1.2150 0.4125 ;
        RECT 1.0500 0.3375 1.1250 0.8250 ;
        RECT 0.7725 0.1650 0.8475 0.8925 ;
        RECT 0.5325 0.1650 0.7725 0.2400 ;
        RECT 0.6825 0.8175 0.7725 0.8925 ;
    END
END XOR3_1010


MACRO XOR4_0011
    CLASS CORE ;
    FOREIGN XOR4_0011 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.4100 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 2.8200 0.7125 3.2850 0.7875 ;
        RECT 2.8200 0.2625 2.9625 0.3375 ;
        RECT 2.7450 0.2625 2.8200 0.7875 ;
        VIA 2.8800 0.7500 VIA12_square ;
        VIA 2.8500 0.3000 VIA12_square ;
        END
    END Z
    PIN A4
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.5175 0.5625 0.7125 0.6375 ;
        RECT 0.3525 0.4950 0.5175 0.6375 ;
        RECT 0.1725 0.5625 0.3525 0.6375 ;
        VIA 0.4350 0.5400 VIA12_square ;
        END
    END A4
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.3500 0.8625 1.6800 0.9375 ;
        RECT 1.2750 0.5925 1.3500 0.9375 ;
        RECT 1.1400 0.8625 1.2750 0.9375 ;
        VIA 1.3125 0.6750 VIA12_square ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 3.1575 0.4125 3.2775 0.4875 ;
        RECT 3.0825 0.1125 3.1575 0.4875 ;
        RECT 2.5950 0.1125 3.0825 0.1875 ;
        VIA 3.1650 0.4500 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 4.0575 0.5625 4.3200 0.6375 ;
        RECT 3.8925 0.4950 4.0575 0.6375 ;
        RECT 3.7800 0.5625 3.8925 0.6375 ;
        VIA 3.9750 0.5400 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 4.1550 -0.0750 4.4100 0.0750 ;
        RECT 4.0350 -0.0750 4.1550 0.1800 ;
        RECT 3.1200 -0.0750 4.0350 0.0750 ;
        RECT 3.0150 -0.0750 3.1200 0.2550 ;
        RECT 2.7000 -0.0750 3.0150 0.0750 ;
        RECT 2.5950 -0.0750 2.7000 0.2175 ;
        RECT 1.4100 -0.0750 2.5950 0.0750 ;
        RECT 1.3200 -0.0750 1.4100 0.2400 ;
        RECT 0.3750 -0.0750 1.3200 0.0750 ;
        RECT 0.2550 -0.0750 0.3750 0.1875 ;
        RECT 0.0000 -0.0750 0.2550 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 4.1550 0.9750 4.4100 1.1250 ;
        RECT 4.0350 0.8550 4.1550 1.1250 ;
        RECT 3.1050 0.9750 4.0350 1.1250 ;
        RECT 2.9850 0.8625 3.1050 1.1250 ;
        RECT 2.6850 0.9750 2.9850 1.1250 ;
        RECT 2.5650 0.8700 2.6850 1.1250 ;
        RECT 1.4250 0.9750 2.5650 1.1250 ;
        RECT 1.3050 0.8625 1.4250 1.1250 ;
        RECT 0.3750 0.9750 1.3050 1.1250 ;
        RECT 0.2550 0.8625 0.3750 1.1250 ;
        RECT 0.0000 0.9750 0.2550 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 4.2750 0.2700 4.3350 0.3300 ;
        RECT 4.2750 0.8175 4.3350 0.8775 ;
        RECT 4.1625 0.4725 4.2225 0.5325 ;
        RECT 4.0650 0.1200 4.1250 0.1800 ;
        RECT 4.0650 0.8625 4.1250 0.9225 ;
        RECT 3.9675 0.4200 4.0275 0.4800 ;
        RECT 3.9600 0.6600 4.0200 0.7200 ;
        RECT 3.7500 0.6525 3.8100 0.7125 ;
        RECT 3.6450 0.1650 3.7050 0.2250 ;
        RECT 3.6450 0.8325 3.7050 0.8925 ;
        RECT 3.5475 0.3525 3.6075 0.4125 ;
        RECT 3.4350 0.1725 3.4950 0.2325 ;
        RECT 3.4350 0.8325 3.4950 0.8925 ;
        RECT 3.3300 0.4725 3.3900 0.5325 ;
        RECT 3.2250 0.1800 3.2850 0.2400 ;
        RECT 3.2250 0.7200 3.2850 0.7800 ;
        RECT 3.1200 0.5100 3.1800 0.5700 ;
        RECT 3.0150 0.1650 3.0750 0.2250 ;
        RECT 3.0150 0.8625 3.0750 0.9225 ;
        RECT 2.9100 0.4800 2.9700 0.5400 ;
        RECT 2.8050 0.2025 2.8650 0.2625 ;
        RECT 2.8050 0.7200 2.8650 0.7800 ;
        RECT 2.7075 0.4800 2.7675 0.5400 ;
        RECT 2.5950 0.1275 2.6550 0.1875 ;
        RECT 2.5950 0.8700 2.6550 0.9300 ;
        RECT 2.4900 0.4125 2.5500 0.4725 ;
        RECT 2.3850 0.1800 2.4450 0.2400 ;
        RECT 2.2725 0.5850 2.3325 0.6450 ;
        RECT 2.1750 0.2475 2.2350 0.3075 ;
        RECT 2.1750 0.8175 2.2350 0.8775 ;
        RECT 2.0775 0.5850 2.1375 0.6450 ;
        RECT 1.9650 0.2475 2.0250 0.3075 ;
        RECT 1.9650 0.8100 2.0250 0.8700 ;
        RECT 1.8525 0.5400 1.9125 0.6000 ;
        RECT 1.7550 0.2400 1.8150 0.3000 ;
        RECT 1.7550 0.8025 1.8150 0.8625 ;
        RECT 1.5450 0.1725 1.6050 0.2325 ;
        RECT 1.5450 0.7500 1.6050 0.8100 ;
        RECT 1.4400 0.4950 1.5000 0.5550 ;
        RECT 1.3350 0.1500 1.3950 0.2100 ;
        RECT 1.3350 0.8700 1.3950 0.9300 ;
        RECT 1.2300 0.4950 1.2900 0.5550 ;
        RECT 1.1250 0.1800 1.1850 0.2400 ;
        RECT 1.1250 0.7200 1.1850 0.7800 ;
        RECT 1.0200 0.4950 1.0800 0.5550 ;
        RECT 0.9150 0.1725 0.9750 0.2325 ;
        RECT 0.9150 0.8325 0.9750 0.8925 ;
        RECT 0.8100 0.3525 0.8700 0.4125 ;
        RECT 0.7050 0.1650 0.7650 0.2250 ;
        RECT 0.7050 0.8325 0.7650 0.8925 ;
        RECT 0.6000 0.6525 0.6600 0.7125 ;
        RECT 0.3900 0.6600 0.4500 0.7200 ;
        RECT 0.3825 0.4200 0.4425 0.4800 ;
        RECT 0.2850 0.1200 0.3450 0.1800 ;
        RECT 0.2850 0.8700 0.3450 0.9300 ;
        RECT 0.1875 0.4725 0.2475 0.5325 ;
        RECT 0.0750 0.2700 0.1350 0.3300 ;
        RECT 0.0750 0.8175 0.1350 0.8775 ;
        LAYER M1 ;
        RECT 4.2975 0.2625 4.3725 0.9000 ;
        RECT 4.1100 0.2625 4.2975 0.3375 ;
        RECT 4.2525 0.6900 4.2975 0.9000 ;
        RECT 4.0500 0.6900 4.2525 0.7650 ;
        RECT 4.0425 0.4425 4.2225 0.5775 ;
        RECT 3.9300 0.6600 4.0500 0.7650 ;
        RECT 3.9675 0.3900 4.0425 0.5775 ;
        RECT 3.8925 0.4875 3.9675 0.5775 ;
        RECT 3.7275 0.1500 3.9300 0.2325 ;
        RECT 3.7875 0.3075 3.8925 0.4125 ;
        RECT 3.4125 0.4875 3.8925 0.5625 ;
        RECT 3.4050 0.8175 3.8550 0.9000 ;
        RECT 3.7200 0.6375 3.8400 0.7425 ;
        RECT 3.5175 0.3300 3.7875 0.4125 ;
        RECT 3.5925 0.1500 3.7275 0.2550 ;
        RECT 3.2925 0.6675 3.7200 0.7425 ;
        RECT 3.3600 0.1500 3.5175 0.2550 ;
        RECT 3.3000 0.4425 3.4125 0.5625 ;
        RECT 3.2100 0.1500 3.3600 0.3000 ;
        RECT 3.2175 0.6675 3.2925 0.8100 ;
        RECT 3.0525 0.3750 3.2175 0.5925 ;
        RECT 2.8575 0.6675 3.0300 0.7875 ;
        RECT 2.7825 0.4500 2.9700 0.5700 ;
        RECT 2.7750 0.1500 2.9400 0.3750 ;
        RECT 2.5875 0.7125 2.8575 0.7875 ;
        RECT 2.7075 0.4500 2.7825 0.6375 ;
        RECT 2.4825 0.5625 2.7075 0.6375 ;
        RECT 2.5575 0.3225 2.6325 0.4875 ;
        RECT 2.4375 0.4050 2.5575 0.4875 ;
        RECT 2.4825 0.1500 2.5200 0.2550 ;
        RECT 2.3100 0.1500 2.4825 0.3300 ;
        RECT 2.4075 0.5625 2.4825 0.9000 ;
        RECT 2.2350 0.4050 2.4375 0.4800 ;
        RECT 1.9650 0.7800 2.4075 0.9000 ;
        RECT 1.9875 0.5550 2.3325 0.6900 ;
        RECT 2.1450 0.1950 2.2350 0.4800 ;
        RECT 1.9350 0.1950 2.0700 0.4350 ;
        RECT 1.8075 0.5100 1.9125 0.6300 ;
        RECT 1.7250 0.7050 1.8900 0.9000 ;
        RECT 1.7475 0.1500 1.8600 0.4350 ;
        RECT 1.6500 0.5100 1.8075 0.5850 ;
        RECT 1.5750 0.1500 1.6500 0.8175 ;
        RECT 1.5075 0.1500 1.5750 0.2550 ;
        RECT 1.5150 0.7425 1.5750 0.8175 ;
        RECT 1.4250 0.3300 1.5000 0.6375 ;
        RECT 1.3200 0.3300 1.4250 0.4125 ;
        RECT 1.2600 0.4875 1.3500 0.7575 ;
        RECT 1.1850 0.4875 1.2600 0.5925 ;
        RECT 1.0425 0.1500 1.2000 0.4125 ;
        RECT 1.1100 0.6675 1.1850 0.8100 ;
        RECT 1.0050 0.4875 1.1100 0.5925 ;
        RECT 0.6900 0.6675 1.1100 0.7425 ;
        RECT 0.8925 0.1500 1.0425 0.2550 ;
        RECT 0.5175 0.4875 1.0050 0.5625 ;
        RECT 0.5550 0.8175 1.0050 0.9000 ;
        RECT 0.6225 0.3300 0.9375 0.4125 ;
        RECT 0.7125 0.1500 0.8175 0.2550 ;
        RECT 0.4800 0.1500 0.7125 0.2325 ;
        RECT 0.5700 0.6375 0.6900 0.7425 ;
        RECT 0.5175 0.3075 0.6225 0.4125 ;
        RECT 0.4425 0.4875 0.5175 0.5775 ;
        RECT 0.1575 0.6600 0.4800 0.7650 ;
        RECT 0.3450 0.3900 0.4425 0.5775 ;
        RECT 0.1875 0.4425 0.3450 0.5775 ;
        RECT 0.1125 0.2625 0.2850 0.3375 ;
        RECT 0.1125 0.6600 0.1575 0.9000 ;
        RECT 0.0375 0.2625 0.1125 0.9000 ;
        LAYER VIA1 ;
        RECT 4.1550 0.2625 4.2300 0.3375 ;
        RECT 3.7725 0.3300 3.8475 0.4050 ;
        RECT 3.6375 0.1575 3.7125 0.2325 ;
        RECT 3.5850 0.8175 3.6600 0.8925 ;
        RECT 3.4350 0.6675 3.5100 0.7425 ;
        RECT 3.3900 0.1650 3.4650 0.2400 ;
        RECT 2.5125 0.4125 2.5875 0.4875 ;
        RECT 2.4075 0.6975 2.4825 0.7725 ;
        RECT 2.3550 0.1725 2.4300 0.2475 ;
        RECT 2.0325 0.5775 2.1075 0.6525 ;
        RECT 1.9650 0.3300 2.0400 0.4050 ;
        RECT 1.8150 0.7800 1.8900 0.8550 ;
        RECT 1.7700 0.2100 1.8450 0.2850 ;
        RECT 1.3800 0.3375 1.4550 0.4125 ;
        RECT 1.0875 0.3225 1.1625 0.3975 ;
        RECT 1.0425 0.6675 1.1175 0.7425 ;
        RECT 0.8250 0.8175 0.9000 0.8925 ;
        RECT 0.6975 0.1575 0.7725 0.2325 ;
        RECT 0.5625 0.3375 0.6375 0.4125 ;
        RECT 0.1650 0.2625 0.2400 0.3375 ;
        LAYER M2 ;
        RECT 4.0200 0.2625 4.2750 0.3375 ;
        RECT 3.9450 0.2625 4.0200 0.4200 ;
        RECT 3.7350 0.3150 3.9450 0.4200 ;
        RECT 3.6600 0.1575 3.7875 0.2325 ;
        RECT 3.5850 0.1575 3.6600 0.9375 ;
        RECT 2.6700 0.8625 3.5850 0.9375 ;
        RECT 3.4350 0.1500 3.5100 0.7875 ;
        RECT 3.3525 0.1500 3.4350 0.2550 ;
        RECT 3.4050 0.6825 3.4350 0.7875 ;
        RECT 2.5950 0.4125 2.6700 0.9375 ;
        RECT 2.4675 0.4125 2.5950 0.4875 ;
        RECT 1.9050 0.8625 2.5950 0.9375 ;
        RECT 2.3025 0.6825 2.5200 0.7875 ;
        RECT 2.3100 0.1650 2.4750 0.2625 ;
        RECT 1.8525 0.1650 2.3100 0.2400 ;
        RECT 2.2275 0.3450 2.3025 0.7875 ;
        RECT 2.0775 0.3450 2.2275 0.4200 ;
        RECT 1.9875 0.5625 2.1525 0.6675 ;
        RECT 1.9275 0.3150 2.0775 0.4200 ;
        RECT 1.5900 0.5625 1.9875 0.6375 ;
        RECT 1.8000 0.7350 1.9050 0.9375 ;
        RECT 1.7475 0.1650 1.8525 0.3300 ;
        RECT 1.5150 0.3375 1.5900 0.6375 ;
        RECT 1.4175 0.3375 1.5150 0.4125 ;
        RECT 1.3350 0.1575 1.4175 0.4125 ;
        RECT 0.9525 0.1575 1.3350 0.2325 ;
        RECT 1.1325 0.3150 1.2075 0.4200 ;
        RECT 1.0275 0.3150 1.1325 0.7875 ;
        RECT 0.8775 0.1575 0.9525 0.9000 ;
        RECT 0.6525 0.1575 0.8775 0.2325 ;
        RECT 0.7800 0.7950 0.8775 0.9000 ;
        RECT 0.5100 0.3375 0.6825 0.4125 ;
        RECT 0.4350 0.2625 0.5100 0.4125 ;
        RECT 0.1200 0.2625 0.4350 0.3375 ;
    END
END XOR4_0011


MACRO XOR4_0111
    CLASS CORE ;
    FOREIGN XOR4_0111 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.3000 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 3.3075 0.2625 3.6225 0.7125 ;
        VIA 3.4650 0.3225 VIA12_slot ;
        VIA 3.4650 0.6525 VIA12_slot ;
        END
    END Z
    PIN A4
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.5175 0.5625 0.7125 0.6375 ;
        RECT 0.3525 0.4950 0.5175 0.6375 ;
        RECT 0.1725 0.5625 0.3525 0.6375 ;
        VIA 0.4350 0.5400 VIA12_square ;
        END
    END A4
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.3500 0.8625 1.6125 0.9375 ;
        RECT 1.2750 0.5925 1.3500 0.9375 ;
        RECT 1.0725 0.8625 1.2750 0.9375 ;
        VIA 1.3125 0.6750 VIA12_square ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 4.1475 0.4125 4.2975 0.4875 ;
        RECT 4.0425 0.4125 4.1475 0.6075 ;
        RECT 3.7575 0.4125 4.0425 0.4875 ;
        VIA 4.0950 0.5250 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 5.3400 0.4125 6.1575 0.4875 ;
        RECT 5.2650 0.3225 5.3400 0.4875 ;
        RECT 4.7025 0.3225 5.2650 0.4050 ;
        RECT 4.6275 0.3225 4.7025 0.4950 ;
        VIA 6.0450 0.4500 VIA12_square ;
        VIA 5.3925 0.4500 VIA12_square ;
        VIA 4.6650 0.4125 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 6.2475 -0.0750 6.3000 0.0750 ;
        RECT 6.1425 -0.0750 6.2475 0.2700 ;
        RECT 5.4150 -0.0750 6.1425 0.0750 ;
        RECT 5.2950 -0.0750 5.4150 0.1875 ;
        RECT 4.3425 -0.0750 5.2950 0.0750 ;
        RECT 4.2375 -0.0750 4.3425 0.2475 ;
        RECT 3.9225 -0.0750 4.2375 0.0750 ;
        RECT 3.8475 -0.0750 3.9225 0.3150 ;
        RECT 3.5250 -0.0750 3.8475 0.0750 ;
        RECT 3.4050 -0.0750 3.5250 0.2025 ;
        RECT 3.0900 -0.0750 3.4050 0.0750 ;
        RECT 3.0150 -0.0750 3.0900 0.2625 ;
        RECT 2.6550 -0.0750 3.0150 0.0750 ;
        RECT 2.5800 -0.0750 2.6550 0.2625 ;
        RECT 1.4100 -0.0750 2.5800 0.0750 ;
        RECT 1.3200 -0.0750 1.4100 0.2400 ;
        RECT 0.3750 -0.0750 1.3200 0.0750 ;
        RECT 0.2550 -0.0750 0.3750 0.1875 ;
        RECT 0.0000 -0.0750 0.2550 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 6.0450 0.9750 6.3000 1.1250 ;
        RECT 5.9400 0.8100 6.0450 1.1250 ;
        RECT 5.6175 0.9750 5.9400 1.1250 ;
        RECT 5.5125 0.7875 5.6175 1.1250 ;
        RECT 4.3650 0.9750 5.5125 1.1250 ;
        RECT 4.2450 0.8025 4.3650 1.1250 ;
        RECT 3.9450 0.9750 4.2450 1.1250 ;
        RECT 3.8250 0.6525 3.9450 1.1250 ;
        RECT 3.5100 0.9750 3.8250 1.1250 ;
        RECT 3.4200 0.8025 3.5100 1.1250 ;
        RECT 3.0900 0.9750 3.4200 1.1250 ;
        RECT 3.0000 0.7650 3.0900 1.1250 ;
        RECT 2.6850 0.9750 3.0000 1.1250 ;
        RECT 2.5650 0.8700 2.6850 1.1250 ;
        RECT 1.4250 0.9750 2.5650 1.1250 ;
        RECT 1.3050 0.8625 1.4250 1.1250 ;
        RECT 0.3750 0.9750 1.3050 1.1250 ;
        RECT 0.2550 0.8625 0.3750 1.1250 ;
        RECT 0.0000 0.9750 0.2550 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 6.1650 0.1875 6.2250 0.2475 ;
        RECT 6.1650 0.6900 6.2250 0.7500 ;
        RECT 6.0600 0.4725 6.1200 0.5325 ;
        RECT 5.9550 0.1725 6.0150 0.2325 ;
        RECT 5.9550 0.8400 6.0150 0.9000 ;
        RECT 5.8500 0.4800 5.9100 0.5400 ;
        RECT 5.7450 0.8175 5.8050 0.8775 ;
        RECT 5.6400 0.4800 5.7000 0.5400 ;
        RECT 5.5350 0.2700 5.5950 0.3300 ;
        RECT 5.5350 0.8175 5.5950 0.8775 ;
        RECT 5.4300 0.4650 5.4900 0.5250 ;
        RECT 5.3250 0.1200 5.3850 0.1800 ;
        RECT 5.2200 0.4650 5.2800 0.5250 ;
        RECT 5.1150 0.2400 5.1750 0.3000 ;
        RECT 5.1150 0.8175 5.1750 0.8775 ;
        RECT 5.0100 0.6450 5.0700 0.7050 ;
        RECT 4.9050 0.2325 4.9650 0.2925 ;
        RECT 4.9050 0.8175 4.9650 0.8775 ;
        RECT 4.8000 0.4875 4.8600 0.5475 ;
        RECT 4.6950 0.1725 4.7550 0.2325 ;
        RECT 4.6950 0.8250 4.7550 0.8850 ;
        RECT 4.5900 0.4500 4.6500 0.5100 ;
        RECT 4.4850 0.6525 4.5450 0.7125 ;
        RECT 4.2750 0.1575 4.3350 0.2175 ;
        RECT 4.2750 0.8100 4.3350 0.8700 ;
        RECT 4.1700 0.4875 4.2300 0.5475 ;
        RECT 4.0650 0.3075 4.1250 0.3675 ;
        RECT 4.0650 0.7275 4.1250 0.7875 ;
        RECT 3.9600 0.4875 4.0200 0.5475 ;
        RECT 3.8550 0.2250 3.9150 0.2850 ;
        RECT 3.8550 0.6675 3.9150 0.7275 ;
        RECT 3.8550 0.8325 3.9150 0.8925 ;
        RECT 3.7500 0.4650 3.8100 0.5250 ;
        RECT 3.6450 0.2250 3.7050 0.2850 ;
        RECT 3.6450 0.7575 3.7050 0.8175 ;
        RECT 3.5400 0.4650 3.6000 0.5250 ;
        RECT 3.4350 0.1350 3.4950 0.1950 ;
        RECT 3.4350 0.8325 3.4950 0.8925 ;
        RECT 3.3300 0.4650 3.3900 0.5250 ;
        RECT 3.2250 0.2250 3.2850 0.2850 ;
        RECT 3.2250 0.7575 3.2850 0.8175 ;
        RECT 3.1200 0.4650 3.1800 0.5250 ;
        RECT 3.0150 0.1725 3.0750 0.2325 ;
        RECT 3.0150 0.8025 3.0750 0.8625 ;
        RECT 2.9100 0.3975 2.9700 0.4575 ;
        RECT 2.8050 0.1725 2.8650 0.2325 ;
        RECT 2.8050 0.7275 2.8650 0.7875 ;
        RECT 2.7000 0.4125 2.7600 0.4725 ;
        RECT 2.5950 0.1725 2.6550 0.2325 ;
        RECT 2.5950 0.8700 2.6550 0.9300 ;
        RECT 2.4900 0.4125 2.5500 0.4725 ;
        RECT 2.3850 0.7800 2.4450 0.8400 ;
        RECT 2.1750 0.2175 2.2350 0.2775 ;
        RECT 2.1750 0.8250 2.2350 0.8850 ;
        RECT 2.0700 0.5025 2.1300 0.5625 ;
        RECT 1.9650 0.2400 2.0250 0.3000 ;
        RECT 1.9650 0.7200 2.0250 0.7800 ;
        RECT 1.8600 0.5025 1.9200 0.5625 ;
        RECT 1.7550 0.2400 1.8150 0.3000 ;
        RECT 1.7550 0.8100 1.8150 0.8700 ;
        RECT 1.5450 0.1725 1.6050 0.2325 ;
        RECT 1.5450 0.7500 1.6050 0.8100 ;
        RECT 1.4400 0.4950 1.5000 0.5550 ;
        RECT 1.3350 0.1500 1.3950 0.2100 ;
        RECT 1.3350 0.8700 1.3950 0.9300 ;
        RECT 1.2300 0.4950 1.2900 0.5550 ;
        RECT 1.1250 0.1800 1.1850 0.2400 ;
        RECT 1.1250 0.7200 1.1850 0.7800 ;
        RECT 1.0200 0.4950 1.0800 0.5550 ;
        RECT 0.9150 0.1725 0.9750 0.2325 ;
        RECT 0.9150 0.8325 0.9750 0.8925 ;
        RECT 0.8100 0.3525 0.8700 0.4125 ;
        RECT 0.7050 0.1650 0.7650 0.2250 ;
        RECT 0.7050 0.8325 0.7650 0.8925 ;
        RECT 0.6000 0.6525 0.6600 0.7125 ;
        RECT 0.3900 0.6600 0.4500 0.7200 ;
        RECT 0.3825 0.4200 0.4425 0.4800 ;
        RECT 0.2850 0.1200 0.3450 0.1800 ;
        RECT 0.2850 0.8700 0.3450 0.9300 ;
        RECT 0.1875 0.4725 0.2475 0.5325 ;
        RECT 0.0750 0.2700 0.1350 0.3300 ;
        RECT 0.0750 0.8175 0.1350 0.8775 ;
        LAYER M1 ;
        RECT 6.0975 0.4350 6.2550 0.5550 ;
        RECT 6.1500 0.6525 6.2400 0.7875 ;
        RECT 5.9175 0.6525 6.1500 0.7275 ;
        RECT 5.9925 0.3300 6.0975 0.5550 ;
        RECT 5.9175 0.1500 6.0375 0.2550 ;
        RECT 5.8425 0.1500 5.9175 0.7275 ;
        RECT 5.6100 0.4575 5.8425 0.5550 ;
        RECT 5.7675 0.8025 5.8350 0.9000 ;
        RECT 5.6925 0.6375 5.7675 0.9000 ;
        RECT 5.2875 0.6375 5.6925 0.7125 ;
        RECT 5.1825 0.2625 5.6475 0.3375 ;
        RECT 5.1975 0.4125 5.5125 0.5550 ;
        RECT 5.2125 0.6375 5.2875 0.9000 ;
        RECT 5.0925 0.7950 5.2125 0.9000 ;
        RECT 5.1075 0.1950 5.1825 0.3375 ;
        RECT 4.4925 0.6450 5.1075 0.7200 ;
        RECT 4.7775 0.4650 5.0925 0.5700 ;
        RECT 4.8750 0.1500 5.0325 0.3600 ;
        RECT 4.6425 0.7950 4.9875 0.9000 ;
        RECT 4.4925 0.1500 4.7775 0.2550 ;
        RECT 4.5675 0.3300 4.7025 0.5700 ;
        RECT 4.4175 0.1500 4.4925 0.7200 ;
        RECT 4.1550 0.3225 4.4175 0.3975 ;
        RECT 4.1325 0.6450 4.4175 0.7200 ;
        RECT 4.0425 0.4800 4.3050 0.5700 ;
        RECT 4.1100 0.2775 4.1550 0.3975 ;
        RECT 4.0575 0.6450 4.1325 0.8250 ;
        RECT 4.0350 0.2775 4.1100 0.3900 ;
        RECT 3.9375 0.4650 4.0425 0.5700 ;
        RECT 3.7500 0.4425 3.8400 0.5400 ;
        RECT 3.1425 0.4425 3.7500 0.5325 ;
        RECT 3.6225 0.1950 3.7275 0.3675 ;
        RECT 3.6375 0.6075 3.7125 0.8700 ;
        RECT 3.2925 0.6075 3.6375 0.6975 ;
        RECT 3.3075 0.2775 3.6225 0.3675 ;
        RECT 3.2025 0.1950 3.3075 0.3675 ;
        RECT 3.2175 0.6075 3.2925 0.8700 ;
        RECT 3.0675 0.4425 3.1425 0.6450 ;
        RECT 2.6400 0.5550 3.0675 0.6450 ;
        RECT 2.8425 0.3750 2.9925 0.4800 ;
        RECT 2.7300 0.1500 2.9400 0.3000 ;
        RECT 2.4525 0.7200 2.8950 0.7950 ;
        RECT 2.4600 0.4050 2.8425 0.4800 ;
        RECT 2.3850 0.1875 2.4600 0.4800 ;
        RECT 2.3775 0.7200 2.4525 0.8925 ;
        RECT 2.1750 0.1875 2.3850 0.3075 ;
        RECT 2.1450 0.8175 2.3775 0.8925 ;
        RECT 2.0175 0.4650 2.3100 0.5850 ;
        RECT 2.0400 0.6600 2.2650 0.7425 ;
        RECT 1.9350 0.1500 2.1000 0.3900 ;
        RECT 1.9500 0.6600 2.0400 0.8250 ;
        RECT 1.8375 0.4725 1.9425 0.5850 ;
        RECT 1.7325 0.6600 1.8675 0.9000 ;
        RECT 1.7325 0.1500 1.8600 0.3975 ;
        RECT 1.6500 0.5100 1.8375 0.5850 ;
        RECT 1.5750 0.1500 1.6500 0.8175 ;
        RECT 1.5075 0.1500 1.5750 0.2550 ;
        RECT 1.5150 0.7425 1.5750 0.8175 ;
        RECT 1.4250 0.3300 1.5000 0.6375 ;
        RECT 1.3200 0.3300 1.4250 0.4125 ;
        RECT 1.2600 0.4875 1.3500 0.7575 ;
        RECT 1.1850 0.4875 1.2600 0.5925 ;
        RECT 1.0425 0.1500 1.2000 0.4125 ;
        RECT 1.1100 0.6675 1.1850 0.8100 ;
        RECT 1.0050 0.4875 1.1100 0.5925 ;
        RECT 0.6900 0.6675 1.1100 0.7425 ;
        RECT 0.8925 0.1500 1.0425 0.2550 ;
        RECT 0.5175 0.4875 1.0050 0.5625 ;
        RECT 0.5550 0.8175 1.0050 0.9000 ;
        RECT 0.6225 0.3300 0.9375 0.4125 ;
        RECT 0.7125 0.1500 0.8175 0.2550 ;
        RECT 0.4800 0.1500 0.7125 0.2325 ;
        RECT 0.5700 0.6375 0.6900 0.7425 ;
        RECT 0.5175 0.3075 0.6225 0.4125 ;
        RECT 0.4425 0.4875 0.5175 0.5775 ;
        RECT 0.1575 0.6600 0.4800 0.7650 ;
        RECT 0.3450 0.3900 0.4425 0.5775 ;
        RECT 0.1875 0.4425 0.3450 0.5775 ;
        RECT 0.1125 0.2625 0.2850 0.3375 ;
        RECT 0.1125 0.6600 0.1575 0.9000 ;
        RECT 0.0375 0.2625 0.1125 0.9000 ;
        LAYER VIA1 ;
        RECT 5.8425 0.6075 5.9175 0.6825 ;
        RECT 4.9500 0.4950 5.0250 0.5700 ;
        RECT 4.9125 0.1650 4.9875 0.2400 ;
        RECT 4.7625 0.8100 4.8375 0.8850 ;
        RECT 2.8800 0.3900 2.9550 0.4650 ;
        RECT 2.7900 0.1650 2.8650 0.2400 ;
        RECT 2.6850 0.5625 2.7600 0.6375 ;
        RECT 2.1750 0.4650 2.2500 0.5400 ;
        RECT 2.0475 0.6600 2.1225 0.7350 ;
        RECT 1.9800 0.3150 2.0550 0.3900 ;
        RECT 1.7625 0.7725 1.8375 0.8475 ;
        RECT 1.7475 0.2100 1.8225 0.2850 ;
        RECT 1.3800 0.3375 1.4550 0.4125 ;
        RECT 1.0875 0.3225 1.1625 0.3975 ;
        RECT 1.0425 0.6675 1.1175 0.7425 ;
        RECT 0.8250 0.8175 0.9000 0.8925 ;
        RECT 0.6975 0.1575 0.7725 0.2325 ;
        RECT 0.5625 0.3375 0.6375 0.4125 ;
        RECT 0.1650 0.2625 0.2400 0.3375 ;
        LAYER M2 ;
        RECT 5.8275 0.5625 5.9325 0.7275 ;
        RECT 5.1450 0.5625 5.8275 0.6375 ;
        RECT 5.0700 0.4950 5.1450 0.6375 ;
        RECT 4.8975 0.4950 5.0700 0.5700 ;
        RECT 4.5525 0.1650 5.0325 0.2400 ;
        RECT 4.5525 0.8100 4.8825 0.8850 ;
        RECT 4.4775 0.1650 4.5525 0.8850 ;
        RECT 2.9925 0.8100 4.4775 0.8850 ;
        RECT 2.9175 0.3750 2.9925 0.8850 ;
        RECT 2.8425 0.3750 2.9175 0.4800 ;
        RECT 1.8525 0.8100 2.9175 0.8850 ;
        RECT 1.8375 0.1650 2.9100 0.2400 ;
        RECT 2.6850 0.3150 2.7600 0.7350 ;
        RECT 2.0400 0.3150 2.6850 0.3900 ;
        RECT 1.9725 0.6600 2.6850 0.7350 ;
        RECT 2.1600 0.4650 2.3250 0.5400 ;
        RECT 2.1000 0.4650 2.1600 0.5700 ;
        RECT 1.5900 0.4950 2.1000 0.5700 ;
        RECT 1.9350 0.3150 2.0400 0.4200 ;
        RECT 1.7475 0.7350 1.8525 0.8850 ;
        RECT 1.7325 0.1650 1.8375 0.3300 ;
        RECT 1.5150 0.3375 1.5900 0.5700 ;
        RECT 1.4175 0.3375 1.5150 0.4125 ;
        RECT 1.3350 0.1575 1.4175 0.4125 ;
        RECT 0.9525 0.1575 1.3350 0.2325 ;
        RECT 1.1325 0.3150 1.2075 0.4200 ;
        RECT 1.0275 0.3150 1.1325 0.7875 ;
        RECT 0.8775 0.1575 0.9525 0.9000 ;
        RECT 0.6525 0.1575 0.8775 0.2325 ;
        RECT 0.7800 0.7950 0.8775 0.9000 ;
        RECT 0.5100 0.3375 0.6825 0.4125 ;
        RECT 0.4350 0.2625 0.5100 0.4125 ;
        RECT 0.1200 0.2625 0.4350 0.3375 ;
    END
END XOR4_0111


MACRO XOR4_1000
    CLASS CORE ;
    FOREIGN XOR4_1000 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.4100 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 2.3175 0.7125 2.7825 0.7875 ;
        VIA 2.6700 0.7500 VIA12_square ;
        END
    END Z
    PIN A4
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.5175 0.5625 0.7125 0.6375 ;
        RECT 0.3525 0.4950 0.5175 0.6375 ;
        RECT 0.1725 0.5625 0.3525 0.6375 ;
        VIA 0.4350 0.5400 VIA12_square ;
        END
    END A4
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.3500 0.8625 1.6125 0.9375 ;
        RECT 1.2750 0.5925 1.3500 0.9375 ;
        RECT 1.0725 0.8625 1.2750 0.9375 ;
        VIA 1.3125 0.6750 VIA12_square ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 3.0600 0.1125 3.1350 0.5775 ;
        RECT 2.5950 0.1125 3.0600 0.1875 ;
        VIA 3.0975 0.4950 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 4.0575 0.5625 4.2000 0.6375 ;
        RECT 3.9075 0.4875 4.0575 0.6375 ;
        RECT 3.6600 0.5625 3.9075 0.6375 ;
        VIA 3.9825 0.5400 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 4.1550 -0.0750 4.4100 0.0750 ;
        RECT 4.0350 -0.0750 4.1550 0.1800 ;
        RECT 3.1200 -0.0750 4.0350 0.0750 ;
        RECT 3.0150 -0.0750 3.1200 0.2550 ;
        RECT 2.7000 -0.0750 3.0150 0.0750 ;
        RECT 2.5950 -0.0750 2.7000 0.2175 ;
        RECT 1.4100 -0.0750 2.5950 0.0750 ;
        RECT 1.3200 -0.0750 1.4100 0.2400 ;
        RECT 0.3750 -0.0750 1.3200 0.0750 ;
        RECT 0.2550 -0.0750 0.3750 0.1875 ;
        RECT 0.0000 -0.0750 0.2550 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 4.1550 0.9750 4.4100 1.1250 ;
        RECT 4.0350 0.8550 4.1550 1.1250 ;
        RECT 3.1200 0.9750 4.0350 1.1250 ;
        RECT 3.0150 0.8025 3.1200 1.1250 ;
        RECT 2.6850 0.9750 3.0150 1.1250 ;
        RECT 2.5650 0.8700 2.6850 1.1250 ;
        RECT 1.4250 0.9750 2.5650 1.1250 ;
        RECT 1.3050 0.8625 1.4250 1.1250 ;
        RECT 0.3750 0.9750 1.3050 1.1250 ;
        RECT 0.2550 0.8625 0.3750 1.1250 ;
        RECT 0.0000 0.9750 0.2550 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 4.2750 0.1575 4.3350 0.2175 ;
        RECT 4.2750 0.8175 4.3350 0.8775 ;
        RECT 4.1625 0.4725 4.2225 0.5325 ;
        RECT 4.0650 0.1200 4.1250 0.1800 ;
        RECT 4.0650 0.8625 4.1250 0.9225 ;
        RECT 3.9675 0.4200 4.0275 0.4800 ;
        RECT 3.9675 0.6600 4.0275 0.7200 ;
        RECT 3.7425 0.6525 3.8025 0.7125 ;
        RECT 3.6450 0.1575 3.7050 0.2175 ;
        RECT 3.6450 0.8325 3.7050 0.8925 ;
        RECT 3.5400 0.3525 3.6000 0.4125 ;
        RECT 3.4350 0.1725 3.4950 0.2325 ;
        RECT 3.4350 0.8325 3.4950 0.8925 ;
        RECT 3.3300 0.5100 3.3900 0.5700 ;
        RECT 3.2250 0.1575 3.2850 0.2175 ;
        RECT 3.2250 0.7800 3.2850 0.8400 ;
        RECT 3.1200 0.4800 3.1800 0.5400 ;
        RECT 3.0150 0.1575 3.0750 0.2175 ;
        RECT 3.0150 0.8325 3.0750 0.8925 ;
        RECT 2.8050 0.1575 2.8650 0.2175 ;
        RECT 2.8050 0.8175 2.8650 0.8775 ;
        RECT 2.7075 0.4800 2.7675 0.5400 ;
        RECT 2.5950 0.1275 2.6550 0.1875 ;
        RECT 2.5950 0.8700 2.6550 0.9300 ;
        RECT 2.4900 0.4125 2.5500 0.4725 ;
        RECT 2.3850 0.1575 2.4450 0.2175 ;
        RECT 2.2725 0.5850 2.3325 0.6450 ;
        RECT 2.1750 0.1800 2.2350 0.2400 ;
        RECT 2.1750 0.8175 2.2350 0.8775 ;
        RECT 2.0775 0.5850 2.1375 0.6450 ;
        RECT 1.9650 0.1950 2.0250 0.2550 ;
        RECT 1.9650 0.8175 2.0250 0.8775 ;
        RECT 1.8600 0.5175 1.9200 0.5775 ;
        RECT 1.7550 0.1800 1.8150 0.2400 ;
        RECT 1.7550 0.8175 1.8150 0.8775 ;
        RECT 1.5450 0.1575 1.6050 0.2175 ;
        RECT 1.5450 0.8175 1.6050 0.8775 ;
        RECT 1.4400 0.4950 1.5000 0.5550 ;
        RECT 1.3350 0.1500 1.3950 0.2100 ;
        RECT 1.3350 0.8700 1.3950 0.9300 ;
        RECT 1.2300 0.4950 1.2900 0.5550 ;
        RECT 1.1250 0.1575 1.1850 0.2175 ;
        RECT 1.1250 0.7800 1.1850 0.8400 ;
        RECT 1.0200 0.4950 1.0800 0.5550 ;
        RECT 0.9150 0.1725 0.9750 0.2325 ;
        RECT 0.9150 0.8325 0.9750 0.8925 ;
        RECT 0.8100 0.3525 0.8700 0.4125 ;
        RECT 0.7050 0.1650 0.7650 0.2250 ;
        RECT 0.7050 0.8325 0.7650 0.8925 ;
        RECT 0.6000 0.6525 0.6600 0.7125 ;
        RECT 0.3900 0.6600 0.4500 0.7200 ;
        RECT 0.3825 0.4200 0.4425 0.4800 ;
        RECT 0.2850 0.1200 0.3450 0.1800 ;
        RECT 0.2850 0.8700 0.3450 0.9300 ;
        RECT 0.1875 0.4725 0.2475 0.5325 ;
        RECT 0.0750 0.1575 0.1350 0.2175 ;
        RECT 0.0750 0.8175 0.1350 0.8775 ;
        LAYER M1 ;
        RECT 4.2975 0.1500 4.3725 0.9000 ;
        RECT 4.2450 0.1500 4.2975 0.3375 ;
        RECT 4.2525 0.6900 4.2975 0.9000 ;
        RECT 4.0575 0.6900 4.2525 0.7650 ;
        RECT 4.1100 0.2625 4.2450 0.3375 ;
        RECT 4.0425 0.4425 4.2225 0.5775 ;
        RECT 3.9375 0.6600 4.0575 0.7650 ;
        RECT 3.9675 0.3900 4.0425 0.5775 ;
        RECT 3.4200 0.5025 3.9675 0.5775 ;
        RECT 3.5925 0.1500 3.9300 0.2550 ;
        RECT 3.4725 0.3300 3.8625 0.4275 ;
        RECT 3.4050 0.8175 3.8550 0.9000 ;
        RECT 3.7125 0.6525 3.8325 0.7425 ;
        RECT 3.2925 0.6675 3.7125 0.7425 ;
        RECT 3.3375 0.1500 3.5175 0.2550 ;
        RECT 3.4050 0.5025 3.4200 0.5925 ;
        RECT 3.3000 0.4875 3.4050 0.5925 ;
        RECT 3.1950 0.1500 3.3375 0.3225 ;
        RECT 3.2175 0.6675 3.2925 0.8700 ;
        RECT 3.1350 0.3975 3.2175 0.5925 ;
        RECT 3.0525 0.3975 3.1350 0.6825 ;
        RECT 2.8650 0.1500 2.9400 0.8775 ;
        RECT 2.7750 0.1500 2.8650 0.2550 ;
        RECT 2.7750 0.7125 2.8650 0.8775 ;
        RECT 2.7075 0.4350 2.7825 0.6375 ;
        RECT 2.5875 0.7125 2.7750 0.7875 ;
        RECT 2.4825 0.5625 2.7075 0.6375 ;
        RECT 2.5575 0.3225 2.6325 0.4875 ;
        RECT 2.4375 0.4050 2.5575 0.4875 ;
        RECT 2.4825 0.1500 2.5200 0.2550 ;
        RECT 2.3250 0.1500 2.4825 0.3300 ;
        RECT 2.4075 0.5625 2.4825 0.9000 ;
        RECT 2.2500 0.4050 2.4375 0.4800 ;
        RECT 1.9425 0.7800 2.4075 0.9000 ;
        RECT 2.0550 0.5550 2.3325 0.6900 ;
        RECT 2.1450 0.1500 2.2500 0.4800 ;
        RECT 1.9350 0.1500 2.0700 0.4350 ;
        RECT 1.6500 0.5100 1.9500 0.5850 ;
        RECT 1.7250 0.6600 1.8675 0.9000 ;
        RECT 1.7250 0.1500 1.8600 0.3900 ;
        RECT 1.5750 0.1500 1.6500 0.8850 ;
        RECT 1.5075 0.1500 1.5750 0.2550 ;
        RECT 1.5150 0.7800 1.5750 0.8850 ;
        RECT 1.4250 0.3300 1.5000 0.6375 ;
        RECT 1.3200 0.3300 1.4250 0.4125 ;
        RECT 1.2600 0.4875 1.3500 0.7575 ;
        RECT 1.1850 0.4875 1.2600 0.5925 ;
        RECT 1.0425 0.1500 1.2150 0.4125 ;
        RECT 1.1100 0.6675 1.1850 0.8700 ;
        RECT 1.0050 0.4875 1.1100 0.5925 ;
        RECT 0.6900 0.6675 1.1100 0.7425 ;
        RECT 0.8925 0.1500 1.0425 0.2550 ;
        RECT 0.5175 0.4875 1.0050 0.5625 ;
        RECT 0.5550 0.8175 1.0050 0.9000 ;
        RECT 0.6225 0.3300 0.9375 0.4125 ;
        RECT 0.7050 0.1500 0.8175 0.2550 ;
        RECT 0.4800 0.1500 0.7050 0.2325 ;
        RECT 0.5700 0.6375 0.6900 0.7425 ;
        RECT 0.5175 0.3075 0.6225 0.4125 ;
        RECT 0.4425 0.4875 0.5175 0.5775 ;
        RECT 0.1575 0.6600 0.4800 0.7650 ;
        RECT 0.3450 0.3900 0.4425 0.5775 ;
        RECT 0.1875 0.4425 0.3450 0.5775 ;
        RECT 0.1650 0.2625 0.2850 0.3375 ;
        RECT 0.1125 0.1575 0.1650 0.3375 ;
        RECT 0.1125 0.6600 0.1575 0.9000 ;
        RECT 0.0375 0.1575 0.1125 0.9000 ;
        LAYER VIA1 ;
        RECT 4.1550 0.2625 4.2300 0.3375 ;
        RECT 3.7425 0.3525 3.8175 0.4275 ;
        RECT 3.6375 0.1575 3.7125 0.2325 ;
        RECT 3.4650 0.8175 3.5400 0.8925 ;
        RECT 3.2625 0.6675 3.3375 0.7425 ;
        RECT 3.2475 0.1950 3.3225 0.2700 ;
        RECT 2.5575 0.3675 2.6325 0.4425 ;
        RECT 2.4600 0.5625 2.5350 0.6375 ;
        RECT 2.3625 0.1800 2.4375 0.2550 ;
        RECT 2.1000 0.5700 2.1750 0.6450 ;
        RECT 1.9650 0.3300 2.0400 0.4050 ;
        RECT 1.7775 0.7800 1.8525 0.8550 ;
        RECT 1.7700 0.2100 1.8450 0.2850 ;
        RECT 1.3800 0.3375 1.4550 0.4125 ;
        RECT 1.0875 0.3225 1.1625 0.3975 ;
        RECT 1.0425 0.6675 1.1175 0.7425 ;
        RECT 0.8250 0.8175 0.9000 0.8925 ;
        RECT 0.6975 0.1575 0.7725 0.2325 ;
        RECT 0.5625 0.3375 0.6375 0.4125 ;
        RECT 0.1650 0.2625 0.2400 0.3375 ;
        LAYER M2 ;
        RECT 4.0200 0.2625 4.2750 0.3375 ;
        RECT 3.9450 0.2625 4.0200 0.3825 ;
        RECT 3.8325 0.3075 3.9450 0.3825 ;
        RECT 3.7275 0.3075 3.8325 0.4650 ;
        RECT 3.5400 0.1575 3.7875 0.2325 ;
        RECT 3.4650 0.1575 3.5400 0.9375 ;
        RECT 2.9775 0.8625 3.4650 0.9375 ;
        RECT 3.3150 0.1650 3.3900 0.7575 ;
        RECT 3.2175 0.1650 3.3150 0.3000 ;
        RECT 3.2175 0.6525 3.3150 0.7575 ;
        RECT 2.9025 0.3525 2.9775 0.9375 ;
        RECT 2.5125 0.3525 2.9025 0.4575 ;
        RECT 1.8675 0.8625 2.9025 0.9375 ;
        RECT 2.4000 0.5625 2.5800 0.6375 ;
        RECT 2.3175 0.1650 2.4750 0.2700 ;
        RECT 2.3250 0.4125 2.4000 0.6375 ;
        RECT 2.0775 0.4125 2.3250 0.4875 ;
        RECT 1.8525 0.1650 2.3175 0.2400 ;
        RECT 2.0550 0.5625 2.2200 0.6675 ;
        RECT 1.9275 0.3150 2.0775 0.4875 ;
        RECT 1.5900 0.5625 2.0550 0.6375 ;
        RECT 1.7625 0.7350 1.8675 0.9375 ;
        RECT 1.7475 0.1650 1.8525 0.3300 ;
        RECT 1.5150 0.3375 1.5900 0.6375 ;
        RECT 1.4175 0.3375 1.5150 0.4125 ;
        RECT 1.3350 0.1575 1.4175 0.4125 ;
        RECT 0.9525 0.1575 1.3350 0.2325 ;
        RECT 1.1325 0.3150 1.2075 0.4200 ;
        RECT 1.0275 0.3150 1.1325 0.7875 ;
        RECT 0.8775 0.1575 0.9525 0.9000 ;
        RECT 0.6450 0.1575 0.8775 0.2325 ;
        RECT 0.7800 0.7950 0.8775 0.9000 ;
        RECT 0.4950 0.3375 0.6825 0.4125 ;
        RECT 0.4200 0.2625 0.4950 0.4125 ;
        RECT 0.1200 0.2625 0.4200 0.3375 ;
    END
END XOR4_1000


MACRO XOR4_1010
    CLASS CORE ;
    FOREIGN XOR4_1010 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.4100 BY 1.0500 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT 2.3175 0.7125 2.7825 0.7875 ;
        VIA 2.6700 0.7500 VIA12_square ;
        END
    END Z
    PIN A4
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 0.5175 0.5625 0.7125 0.6375 ;
        RECT 0.3525 0.4950 0.5175 0.6375 ;
        RECT 0.1725 0.5625 0.3525 0.6375 ;
        VIA 0.4350 0.5400 VIA12_square ;
        END
    END A4
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 1.3500 0.8625 1.6800 0.9375 ;
        RECT 1.2750 0.5925 1.3500 0.9375 ;
        RECT 1.1400 0.8625 1.2750 0.9375 ;
        VIA 1.3125 0.6750 VIA12_square ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 3.0600 0.1125 3.1350 0.5325 ;
        RECT 2.5950 0.1125 3.0600 0.1875 ;
        VIA 3.0975 0.4500 VIA12_square ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT 4.0575 0.5625 4.3425 0.6375 ;
        RECT 3.8925 0.4950 4.0575 0.6375 ;
        RECT 3.7125 0.5625 3.8925 0.6375 ;
        VIA 3.9750 0.5400 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 4.1550 -0.0750 4.4100 0.0750 ;
        RECT 4.0350 -0.0750 4.1550 0.1800 ;
        RECT 3.1200 -0.0750 4.0350 0.0750 ;
        RECT 3.0150 -0.0750 3.1200 0.2550 ;
        RECT 2.7000 -0.0750 3.0150 0.0750 ;
        RECT 2.5950 -0.0750 2.7000 0.2175 ;
        RECT 1.4100 -0.0750 2.5950 0.0750 ;
        RECT 1.3200 -0.0750 1.4100 0.2400 ;
        RECT 0.3750 -0.0750 1.3200 0.0750 ;
        RECT 0.2550 -0.0750 0.3750 0.1875 ;
        RECT 0.0000 -0.0750 0.2550 0.0750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT 4.1550 0.9750 4.4100 1.1250 ;
        RECT 4.0350 0.8550 4.1550 1.1250 ;
        RECT 3.1200 0.9750 4.0350 1.1250 ;
        RECT 3.0150 0.8025 3.1200 1.1250 ;
        RECT 2.6850 0.9750 3.0150 1.1250 ;
        RECT 2.5650 0.8700 2.6850 1.1250 ;
        RECT 1.4250 0.9750 2.5650 1.1250 ;
        RECT 1.3050 0.8625 1.4250 1.1250 ;
        RECT 0.3750 0.9750 1.3050 1.1250 ;
        RECT 0.2550 0.8625 0.3750 1.1250 ;
        RECT 0.0000 0.9750 0.2550 1.1250 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT 4.2750 0.2700 4.3350 0.3300 ;
        RECT 4.2750 0.8175 4.3350 0.8775 ;
        RECT 4.1625 0.4725 4.2225 0.5325 ;
        RECT 4.0650 0.1200 4.1250 0.1800 ;
        RECT 4.0650 0.8625 4.1250 0.9225 ;
        RECT 3.9675 0.4200 4.0275 0.4800 ;
        RECT 3.9600 0.6600 4.0200 0.7200 ;
        RECT 3.7500 0.6525 3.8100 0.7125 ;
        RECT 3.6450 0.1650 3.7050 0.2250 ;
        RECT 3.6450 0.8325 3.7050 0.8925 ;
        RECT 3.5400 0.3525 3.6000 0.4125 ;
        RECT 3.4350 0.1725 3.4950 0.2325 ;
        RECT 3.4350 0.8325 3.4950 0.8925 ;
        RECT 3.3300 0.4950 3.3900 0.5550 ;
        RECT 3.2250 0.1800 3.2850 0.2400 ;
        RECT 3.2250 0.7200 3.2850 0.7800 ;
        RECT 3.1200 0.5100 3.1800 0.5700 ;
        RECT 3.0150 0.1650 3.0750 0.2250 ;
        RECT 3.0150 0.8325 3.0750 0.8925 ;
        RECT 2.8050 0.2025 2.8650 0.2625 ;
        RECT 2.8050 0.7200 2.8650 0.7800 ;
        RECT 2.7075 0.4800 2.7675 0.5400 ;
        RECT 2.5950 0.1275 2.6550 0.1875 ;
        RECT 2.5950 0.8700 2.6550 0.9300 ;
        RECT 2.4900 0.4125 2.5500 0.4725 ;
        RECT 2.3850 0.1800 2.4450 0.2400 ;
        RECT 2.2725 0.5850 2.3325 0.6450 ;
        RECT 2.1750 0.2475 2.2350 0.3075 ;
        RECT 2.1750 0.8175 2.2350 0.8775 ;
        RECT 2.0775 0.5850 2.1375 0.6450 ;
        RECT 1.9650 0.2475 2.0250 0.3075 ;
        RECT 1.9650 0.8100 2.0250 0.8700 ;
        RECT 1.8600 0.5175 1.9200 0.5775 ;
        RECT 1.7550 0.2400 1.8150 0.3000 ;
        RECT 1.7550 0.8025 1.8150 0.8625 ;
        RECT 1.5450 0.1725 1.6050 0.2325 ;
        RECT 1.5450 0.7500 1.6050 0.8100 ;
        RECT 1.4400 0.4950 1.5000 0.5550 ;
        RECT 1.3350 0.1500 1.3950 0.2100 ;
        RECT 1.3350 0.8700 1.3950 0.9300 ;
        RECT 1.2300 0.4950 1.2900 0.5550 ;
        RECT 1.1250 0.1800 1.1850 0.2400 ;
        RECT 1.1250 0.7200 1.1850 0.7800 ;
        RECT 1.0200 0.4950 1.0800 0.5550 ;
        RECT 0.9150 0.1725 0.9750 0.2325 ;
        RECT 0.9150 0.8325 0.9750 0.8925 ;
        RECT 0.8100 0.3525 0.8700 0.4125 ;
        RECT 0.7050 0.1650 0.7650 0.2250 ;
        RECT 0.7050 0.8325 0.7650 0.8925 ;
        RECT 0.6000 0.6525 0.6600 0.7125 ;
        RECT 0.3900 0.6600 0.4500 0.7200 ;
        RECT 0.3825 0.4200 0.4425 0.4800 ;
        RECT 0.2850 0.1200 0.3450 0.1800 ;
        RECT 0.2850 0.8700 0.3450 0.9300 ;
        RECT 0.1875 0.4725 0.2475 0.5325 ;
        RECT 0.0750 0.2700 0.1350 0.3300 ;
        RECT 0.0750 0.8175 0.1350 0.8775 ;
        LAYER M1 ;
        RECT 4.2975 0.2625 4.3725 0.9000 ;
        RECT 4.1100 0.2625 4.2975 0.3375 ;
        RECT 4.2525 0.6900 4.2975 0.9000 ;
        RECT 4.0500 0.6900 4.2525 0.7650 ;
        RECT 4.0425 0.4425 4.2225 0.5775 ;
        RECT 3.9300 0.6600 4.0500 0.7650 ;
        RECT 3.9675 0.3900 4.0425 0.5775 ;
        RECT 3.8925 0.4875 3.9675 0.5775 ;
        RECT 3.7275 0.1500 3.9300 0.2325 ;
        RECT 3.7875 0.3075 3.8925 0.4125 ;
        RECT 3.4050 0.4875 3.8925 0.5625 ;
        RECT 3.4050 0.8175 3.8550 0.9000 ;
        RECT 3.7200 0.6375 3.8400 0.7425 ;
        RECT 3.4725 0.3300 3.7875 0.4125 ;
        RECT 3.5925 0.1500 3.7275 0.2550 ;
        RECT 3.2925 0.6675 3.7200 0.7425 ;
        RECT 3.3375 0.1500 3.5175 0.2550 ;
        RECT 3.3000 0.4875 3.4050 0.5925 ;
        RECT 3.2100 0.1500 3.3375 0.4050 ;
        RECT 3.2175 0.6675 3.2925 0.8100 ;
        RECT 3.1350 0.4875 3.2175 0.5925 ;
        RECT 3.0525 0.3675 3.1350 0.6825 ;
        RECT 2.8650 0.1725 2.9400 0.7875 ;
        RECT 2.8050 0.1725 2.8650 0.2925 ;
        RECT 2.5875 0.7125 2.8650 0.7875 ;
        RECT 2.7075 0.4350 2.7825 0.6375 ;
        RECT 2.4825 0.5625 2.7075 0.6375 ;
        RECT 2.5575 0.3225 2.6325 0.4875 ;
        RECT 2.4375 0.4050 2.5575 0.4875 ;
        RECT 2.4825 0.1500 2.5200 0.2550 ;
        RECT 2.3100 0.1500 2.4825 0.3300 ;
        RECT 2.4075 0.5625 2.4825 0.9000 ;
        RECT 2.2350 0.4050 2.4375 0.4800 ;
        RECT 1.9650 0.7800 2.4075 0.9000 ;
        RECT 2.0550 0.5550 2.3325 0.6900 ;
        RECT 2.1450 0.1950 2.2350 0.4800 ;
        RECT 1.9350 0.1950 2.0700 0.4350 ;
        RECT 1.6500 0.5100 1.9500 0.5850 ;
        RECT 1.7550 0.6600 1.8900 0.9000 ;
        RECT 1.7475 0.1500 1.8600 0.4350 ;
        RECT 1.5750 0.1500 1.6500 0.8175 ;
        RECT 1.5075 0.1500 1.5750 0.2550 ;
        RECT 1.5150 0.7425 1.5750 0.8175 ;
        RECT 1.4250 0.3300 1.5000 0.6375 ;
        RECT 1.3200 0.3300 1.4250 0.4125 ;
        RECT 1.2600 0.4875 1.3500 0.7575 ;
        RECT 1.1850 0.4875 1.2600 0.5925 ;
        RECT 1.0425 0.1500 1.2000 0.4125 ;
        RECT 1.1100 0.6675 1.1850 0.8100 ;
        RECT 1.0050 0.4875 1.1100 0.5925 ;
        RECT 0.6900 0.6675 1.1100 0.7425 ;
        RECT 0.8925 0.1500 1.0425 0.2550 ;
        RECT 0.5175 0.4875 1.0050 0.5625 ;
        RECT 0.5550 0.8175 1.0050 0.9000 ;
        RECT 0.6225 0.3300 0.9375 0.4125 ;
        RECT 0.7125 0.1500 0.8175 0.2550 ;
        RECT 0.4800 0.1500 0.7125 0.2325 ;
        RECT 0.5700 0.6375 0.6900 0.7425 ;
        RECT 0.5175 0.3075 0.6225 0.4125 ;
        RECT 0.4425 0.4875 0.5175 0.5775 ;
        RECT 0.1575 0.6600 0.4800 0.7650 ;
        RECT 0.3450 0.3900 0.4425 0.5775 ;
        RECT 0.1875 0.4425 0.3450 0.5775 ;
        RECT 0.1125 0.2625 0.2850 0.3375 ;
        RECT 0.1125 0.6600 0.1575 0.9000 ;
        RECT 0.0375 0.2625 0.1125 0.9000 ;
        LAYER VIA1 ;
        RECT 4.1550 0.2625 4.2300 0.3375 ;
        RECT 3.7725 0.3300 3.8475 0.4050 ;
        RECT 3.6375 0.1575 3.7125 0.2325 ;
        RECT 3.4650 0.8175 3.5400 0.8925 ;
        RECT 3.2625 0.6675 3.3375 0.7425 ;
        RECT 3.2475 0.1950 3.3225 0.2700 ;
        RECT 2.5575 0.3675 2.6325 0.4425 ;
        RECT 2.4600 0.5625 2.5350 0.6375 ;
        RECT 2.3550 0.1725 2.4300 0.2475 ;
        RECT 2.1000 0.5700 2.1750 0.6450 ;
        RECT 1.9650 0.3300 2.0400 0.4050 ;
        RECT 1.8150 0.7800 1.8900 0.8550 ;
        RECT 1.7700 0.2100 1.8450 0.2850 ;
        RECT 1.3800 0.3375 1.4550 0.4125 ;
        RECT 1.0875 0.3225 1.1625 0.3975 ;
        RECT 1.0425 0.6675 1.1175 0.7425 ;
        RECT 0.8250 0.8175 0.9000 0.8925 ;
        RECT 0.6975 0.1575 0.7725 0.2325 ;
        RECT 0.5625 0.3375 0.6375 0.4125 ;
        RECT 0.1650 0.2625 0.2400 0.3375 ;
        LAYER M2 ;
        RECT 4.0200 0.2625 4.2750 0.3375 ;
        RECT 3.9450 0.2625 4.0200 0.4050 ;
        RECT 3.7275 0.3300 3.9450 0.4050 ;
        RECT 3.5400 0.1575 3.7575 0.2325 ;
        RECT 3.4650 0.1575 3.5400 0.9375 ;
        RECT 2.9775 0.8625 3.4650 0.9375 ;
        RECT 3.3150 0.1650 3.3900 0.7575 ;
        RECT 3.2175 0.1650 3.3150 0.3000 ;
        RECT 3.2175 0.6525 3.3150 0.7575 ;
        RECT 2.9025 0.3525 2.9775 0.9375 ;
        RECT 2.5125 0.3525 2.9025 0.4575 ;
        RECT 1.9050 0.8625 2.9025 0.9375 ;
        RECT 2.4000 0.5625 2.5800 0.6375 ;
        RECT 2.3100 0.1650 2.4750 0.2625 ;
        RECT 2.3250 0.3450 2.4000 0.6375 ;
        RECT 2.0775 0.3450 2.3250 0.4200 ;
        RECT 1.8525 0.1650 2.3100 0.2400 ;
        RECT 2.0550 0.5625 2.2200 0.6675 ;
        RECT 1.9275 0.3150 2.0775 0.4200 ;
        RECT 1.5900 0.5625 2.0550 0.6375 ;
        RECT 1.8000 0.7350 1.9050 0.9375 ;
        RECT 1.7475 0.1650 1.8525 0.3300 ;
        RECT 1.5150 0.3375 1.5900 0.6375 ;
        RECT 1.4175 0.3375 1.5150 0.4125 ;
        RECT 1.3350 0.1575 1.4175 0.4125 ;
        RECT 0.9525 0.1575 1.3350 0.2325 ;
        RECT 1.1325 0.3150 1.2075 0.4200 ;
        RECT 1.0275 0.3150 1.1325 0.7875 ;
        RECT 0.8775 0.1575 0.9525 0.9000 ;
        RECT 0.6525 0.1575 0.8775 0.2325 ;
        RECT 0.7800 0.7950 0.8775 0.9000 ;
        RECT 0.5100 0.3375 0.6825 0.4125 ;
        RECT 0.4350 0.2625 0.5100 0.4125 ;
        RECT 0.1200 0.2625 0.4350 0.3375 ;
    END
END XOR4_1010


VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO adv_dbg_if
  CLASS BLOCK ;
    SIZE 68.8800 BY 67.2000 ;
  FOREIGN adv_dbg_if 0.000000 0.000000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN tms_pad_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 34.7625 0.0000 34.8375 0.5100 ;
    END
  END tms_pad_i
  PIN tck_pad_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 37.2375 66.7800 37.3125 67.2000 ;
    END
  END tck_pad_i
  PIN trstn_pad_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 68.3700 35.3625 68.8800 35.4375 ;
    END
  END trstn_pad_i
  PIN tdi_pad_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 34.7625 0.0000 34.8375 0.5100 ;
    END
  END tdi_pad_i
  PIN tdo_pad_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 34.9275 0.0000 35.0025 0.4200 ;
    END
  END tdo_pad_o
  PIN tdo_padoe_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 33.8625 66.6900 33.9375 67.2000 ;
    END
  END tdo_padoe_o
  PIN test_mode_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 34.0125 66.6900 34.0875 67.2000 ;
    END
  END test_mode_i
  PIN cpu_clk_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 34.1625 0.0000 34.2375 0.5100 ;
    END
  END cpu_clk_i[0]
  PIN cpu_addr_o[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 57.3975 66.7800 57.4725 67.2000 ;
    END
  END cpu_addr_o[15]
  PIN cpu_addr_o[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 65.7975 66.7800 65.8725 67.2000 ;
    END
  END cpu_addr_o[14]
  PIN cpu_addr_o[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 58.8675 66.7800 58.9425 67.2000 ;
    END
  END cpu_addr_o[13]
  PIN cpu_addr_o[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 68.3700 63.8625 68.8800 63.9375 ;
    END
  END cpu_addr_o[12]
  PIN cpu_addr_o[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 68.3700 62.0625 68.8800 62.1375 ;
    END
  END cpu_addr_o[11]
  PIN cpu_addr_o[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 68.3700 59.6625 68.8800 59.7375 ;
    END
  END cpu_addr_o[10]
  PIN cpu_addr_o[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 68.3700 57.8625 68.8800 57.9375 ;
    END
  END cpu_addr_o[9]
  PIN cpu_addr_o[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 68.3700 53.3625 68.8800 53.4375 ;
    END
  END cpu_addr_o[8]
  PIN cpu_addr_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 68.3700 51.5625 68.8800 51.6375 ;
    END
  END cpu_addr_o[7]
  PIN cpu_addr_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 68.3700 49.1625 68.8800 49.2375 ;
    END
  END cpu_addr_o[6]
  PIN cpu_addr_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 68.3700 47.0625 68.8800 47.1375 ;
    END
  END cpu_addr_o[5]
  PIN cpu_addr_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 68.3700 43.1625 68.8800 43.2375 ;
    END
  END cpu_addr_o[4]
  PIN cpu_addr_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 68.3700 40.7625 68.8800 40.8375 ;
    END
  END cpu_addr_o[3]
  PIN cpu_addr_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 68.3700 34.7625 68.8800 34.8375 ;
    END
  END cpu_addr_o[2]
  PIN cpu_addr_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 66.7575 34.5000 68.8800 35.1000 ;
    END
  END cpu_addr_o[1]
  PIN cpu_addr_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 68.3700 34.4625 68.8800 34.5375 ;
    END
  END cpu_addr_o[0]
  PIN cpu_data_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 14.0625 0.5100 14.1375 ;
    END
  END cpu_data_i[31]
  PIN cpu_data_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 13.1625 0.5100 13.2375 ;
    END
  END cpu_data_i[30]
  PIN cpu_data_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 12.8625 0.5100 12.9375 ;
    END
  END cpu_data_i[29]
  PIN cpu_data_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 13.4625 0.5100 13.5375 ;
    END
  END cpu_data_i[28]
  PIN cpu_data_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 15.2625 0.5100 15.3375 ;
    END
  END cpu_data_i[27]
  PIN cpu_data_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 14.9625 0.5100 15.0375 ;
    END
  END cpu_data_i[26]
  PIN cpu_data_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 15.5625 0.5100 15.6375 ;
    END
  END cpu_data_i[25]
  PIN cpu_data_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 13.7625 0.5100 13.8375 ;
    END
  END cpu_data_i[24]
  PIN cpu_data_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 9.8625 0.5100 9.9375 ;
    END
  END cpu_data_i[23]
  PIN cpu_data_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 7.7625 0.5100 7.8375 ;
    END
  END cpu_data_i[22]
  PIN cpu_data_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9.9375 0.0000 10.0125 0.4200 ;
    END
  END cpu_data_i[21]
  PIN cpu_data_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 4.7625 0.5100 4.8375 ;
    END
  END cpu_data_i[20]
  PIN cpu_data_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 2.6625 0.5100 2.7375 ;
    END
  END cpu_data_i[19]
  PIN cpu_data_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1.4625 0.5100 1.5375 ;
    END
  END cpu_data_i[18]
  PIN cpu_data_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6.5775 0.0000 6.6525 0.4200 ;
    END
  END cpu_data_i[17]
  PIN cpu_data_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10.3575 0.0000 10.4325 0.4200 ;
    END
  END cpu_data_i[16]
  PIN cpu_data_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12.2475 0.0000 12.3225 0.4200 ;
    END
  END cpu_data_i[15]
  PIN cpu_data_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11.8275 0.0000 11.9025 0.4200 ;
    END
  END cpu_data_i[14]
  PIN cpu_data_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18.3375 0.0000 18.4125 0.4200 ;
    END
  END cpu_data_i[13]
  PIN cpu_data_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16.6575 0.0000 16.7325 0.4200 ;
    END
  END cpu_data_i[12]
  PIN cpu_data_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12.6675 0.0000 12.7425 0.4200 ;
    END
  END cpu_data_i[11]
  PIN cpu_data_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13.9275 0.0000 14.0025 0.4200 ;
    END
  END cpu_data_i[10]
  PIN cpu_data_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 19.3875 0.0000 19.4625 0.4200 ;
    END
  END cpu_data_i[9]
  PIN cpu_data_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 19.8075 0.0000 19.8825 0.4200 ;
    END
  END cpu_data_i[8]
  PIN cpu_data_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 21.4875 0.0000 21.5625 0.4200 ;
    END
  END cpu_data_i[7]
  PIN cpu_data_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 23.5875 0.0000 23.6625 0.4200 ;
    END
  END cpu_data_i[6]
  PIN cpu_data_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 24.0075 0.0000 24.0825 0.4200 ;
    END
  END cpu_data_i[5]
  PIN cpu_data_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 21.0675 0.0000 21.1425 0.4200 ;
    END
  END cpu_data_i[4]
  PIN cpu_data_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 22.5375 0.0000 22.6125 0.4200 ;
    END
  END cpu_data_i[3]
  PIN cpu_data_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 21.4125 0.0000 21.4875 0.5100 ;
    END
  END cpu_data_i[2]
  PIN cpu_data_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 28.6275 0.0000 28.7025 0.4200 ;
    END
  END cpu_data_i[1]
  PIN cpu_data_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 32.4075 0.0000 32.4825 0.4200 ;
    END
  END cpu_data_i[0]
  PIN cpu_data_o[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 68.3700 22.1625 68.8800 22.2375 ;
    END
  END cpu_data_o[31]
  PIN cpu_data_o[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 46.8975 0.0000 46.9725 0.4200 ;
    END
  END cpu_data_o[30]
  PIN cpu_data_o[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 68.3700 24.2625 68.8800 24.3375 ;
    END
  END cpu_data_o[29]
  PIN cpu_data_o[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 68.3700 23.9625 68.8800 24.0375 ;
    END
  END cpu_data_o[28]
  PIN cpu_data_o[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 68.3700 28.1625 68.8800 28.2375 ;
    END
  END cpu_data_o[27]
  PIN cpu_data_o[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 68.3700 26.3625 68.8800 26.4375 ;
    END
  END cpu_data_o[26]
  PIN cpu_data_o[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 39.3375 66.7800 39.4125 67.2000 ;
    END
  END cpu_data_o[25]
  PIN cpu_data_o[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 68.3700 28.4625 68.8800 28.5375 ;
    END
  END cpu_data_o[24]
  PIN cpu_data_o[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 68.3700 30.2625 68.8800 30.3375 ;
    END
  END cpu_data_o[23]
  PIN cpu_data_o[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 68.3700 24.2625 68.8800 24.3375 ;
    END
  END cpu_data_o[22]
  PIN cpu_data_o[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 68.3700 34.4625 68.8800 34.5375 ;
    END
  END cpu_data_o[21]
  PIN cpu_data_o[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 68.3700 34.1625 68.8800 34.2375 ;
    END
  END cpu_data_o[20]
  PIN cpu_data_o[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 68.3700 32.3625 68.8800 32.4375 ;
    END
  END cpu_data_o[19]
  PIN cpu_data_o[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 66.7575 32.1000 68.8800 32.7000 ;
    END
  END cpu_data_o[18]
  PIN cpu_data_o[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 68.3700 35.0625 68.8800 35.1375 ;
    END
  END cpu_data_o[17]
  PIN cpu_data_o[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 68.3700 38.9625 68.8800 39.0375 ;
    END
  END cpu_data_o[16]
  PIN cpu_data_o[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 68.3700 36.8625 68.8800 36.9375 ;
    END
  END cpu_data_o[15]
  PIN cpu_data_o[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 68.3700 47.0625 68.8800 47.1375 ;
    END
  END cpu_data_o[14]
  PIN cpu_data_o[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 39.1125 66.6900 39.1875 67.2000 ;
    END
  END cpu_data_o[13]
  PIN cpu_data_o[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 48.7875 66.7800 48.8625 67.2000 ;
    END
  END cpu_data_o[12]
  PIN cpu_data_o[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 68.3700 51.5625 68.8800 51.6375 ;
    END
  END cpu_data_o[11]
  PIN cpu_data_o[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 46.4775 66.7800 46.5525 67.2000 ;
    END
  END cpu_data_o[10]
  PIN cpu_data_o[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 38.2125 66.6900 38.2875 67.2000 ;
    END
  END cpu_data_o[9]
  PIN cpu_data_o[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 47.5275 66.7800 47.6025 67.2000 ;
    END
  END cpu_data_o[8]
  PIN cpu_data_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 68.3700 28.1625 68.8800 28.2375 ;
    END
  END cpu_data_o[7]
  PIN cpu_data_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 49.8375 66.7800 49.9125 67.2000 ;
    END
  END cpu_data_o[6]
  PIN cpu_data_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 42.6975 66.7800 42.7725 67.2000 ;
    END
  END cpu_data_o[5]
  PIN cpu_data_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 48.7125 66.6900 48.7875 67.2000 ;
    END
  END cpu_data_o[4]
  PIN cpu_data_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 52.3575 66.7800 52.4325 67.2000 ;
    END
  END cpu_data_o[3]
  PIN cpu_data_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 50.8875 66.7800 50.9625 67.2000 ;
    END
  END cpu_data_o[2]
  PIN cpu_data_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 40.1775 66.7800 40.2525 67.2000 ;
    END
  END cpu_data_o[1]
  PIN cpu_data_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 44.7975 66.7800 44.8725 67.2000 ;
    END
  END cpu_data_o[0]
  PIN cpu_bp_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 29.0475 0.0000 29.1225 0.4200 ;
    END
  END cpu_bp_i[0]
  PIN cpu_stall_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 28.6125 0.0000 28.6875 0.5100 ;
    END
  END cpu_stall_o[0]
  PIN cpu_stb_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 33.0375 0.0000 33.1125 0.4200 ;
    END
  END cpu_stb_o[0]
  PIN cpu_we_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 33.8625 0.0000 33.9375 0.5100 ;
    END
  END cpu_we_o[0]
  PIN cpu_ack_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 36.3975 0.0000 36.4725 0.4200 ;
    END
  END cpu_ack_i[0]
  PIN cpu_rst_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 47.5125 0.5100 47.5875 ;
    END
  END cpu_rst_o[0]
  PIN axi_aclk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 22.7625 0.5100 22.8375 ;
    END
  END axi_aclk
  PIN axi_aresetn
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 22.4625 0.5100 22.5375 ;
    END
  END axi_aresetn
  PIN axi_master_aw_valid
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 19.7625 0.5100 19.8375 ;
    END
  END axi_master_aw_valid
  PIN axi_master_aw_addr[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 44.6625 0.5100 44.7375 ;
    END
  END axi_master_aw_addr[31]
  PIN axi_master_aw_addr[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 24.5625 66.6900 24.6375 67.2000 ;
    END
  END axi_master_aw_addr[30]
  PIN axi_master_aw_addr[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 30.7125 66.6900 30.7875 67.2000 ;
    END
  END axi_master_aw_addr[29]
  PIN axi_master_aw_addr[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 32.2125 66.6900 32.2875 67.2000 ;
    END
  END axi_master_aw_addr[28]
  PIN axi_master_aw_addr[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 32.2125 0.5100 32.2875 ;
    END
  END axi_master_aw_addr[27]
  PIN axi_master_aw_addr[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 33.1125 0.5100 33.1875 ;
    END
  END axi_master_aw_addr[26]
  PIN axi_master_aw_addr[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 32.8125 0.5100 32.8875 ;
    END
  END axi_master_aw_addr[25]
  PIN axi_master_aw_addr[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 37.3125 0.5100 37.3875 ;
    END
  END axi_master_aw_addr[24]
  PIN axi_master_aw_addr[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 39.5625 0.5100 39.6375 ;
    END
  END axi_master_aw_addr[23]
  PIN axi_master_aw_addr[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 25.6125 66.6900 25.6875 67.2000 ;
    END
  END axi_master_aw_addr[22]
  PIN axi_master_aw_addr[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 34.7625 66.6900 34.8375 67.2000 ;
    END
  END axi_master_aw_addr[21]
  PIN axi_master_aw_addr[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 31.6125 66.6900 31.6875 67.2000 ;
    END
  END axi_master_aw_addr[20]
  PIN axi_master_aw_addr[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 21.1125 66.6900 21.1875 67.2000 ;
    END
  END axi_master_aw_addr[19]
  PIN axi_master_aw_addr[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 31.9125 66.6900 31.9875 67.2000 ;
    END
  END axi_master_aw_addr[18]
  PIN axi_master_aw_addr[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17.6625 66.6900 17.7375 67.2000 ;
    END
  END axi_master_aw_addr[17]
  PIN axi_master_aw_addr[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 21.4125 66.6900 21.4875 67.2000 ;
    END
  END axi_master_aw_addr[16]
  PIN axi_master_aw_addr[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14.9625 66.6900 15.0375 67.2000 ;
    END
  END axi_master_aw_addr[15]
  PIN axi_master_aw_addr[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 20.0625 66.6900 20.1375 67.2000 ;
    END
  END axi_master_aw_addr[14]
  PIN axi_master_aw_addr[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16.9125 66.6900 16.9875 67.2000 ;
    END
  END axi_master_aw_addr[13]
  PIN axi_master_aw_addr[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 25.0125 66.6900 25.0875 67.2000 ;
    END
  END axi_master_aw_addr[12]
  PIN axi_master_aw_addr[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12.7125 66.6900 12.7875 67.2000 ;
    END
  END axi_master_aw_addr[11]
  PIN axi_master_aw_addr[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 28.4625 66.6900 28.5375 67.2000 ;
    END
  END axi_master_aw_addr[10]
  PIN axi_master_aw_addr[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 32.6625 66.6900 32.7375 67.2000 ;
    END
  END axi_master_aw_addr[9]
  PIN axi_master_aw_addr[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 34.3125 66.6900 34.3875 67.2000 ;
    END
  END axi_master_aw_addr[8]
  PIN axi_master_aw_addr[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14.5125 66.6900 14.5875 67.2000 ;
    END
  END axi_master_aw_addr[7]
  PIN axi_master_aw_addr[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 27.7125 66.6900 27.7875 67.2000 ;
    END
  END axi_master_aw_addr[6]
  PIN axi_master_aw_addr[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 19.3125 66.6900 19.3875 67.2000 ;
    END
  END axi_master_aw_addr[5]
  PIN axi_master_aw_addr[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 31.1625 66.6900 31.2375 67.2000 ;
    END
  END axi_master_aw_addr[4]
  PIN axi_master_aw_addr[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 21.8625 66.6900 21.9375 67.2000 ;
    END
  END axi_master_aw_addr[3]
  PIN axi_master_aw_addr[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 34.3125 0.5100 34.3875 ;
    END
  END axi_master_aw_addr[2]
  PIN axi_master_aw_addr[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 23.9625 0.5100 24.0375 ;
    END
  END axi_master_aw_addr[1]
  PIN axi_master_aw_addr[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 26.0625 0.5100 26.1375 ;
    END
  END axi_master_aw_addr[0]
  PIN axi_master_aw_prot[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 47.8125 0.5100 47.8875 ;
    END
  END axi_master_aw_prot[2]
  PIN axi_master_aw_prot[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 48.1125 0.5100 48.1875 ;
    END
  END axi_master_aw_prot[1]
  PIN axi_master_aw_prot[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 48.4125 0.5100 48.4875 ;
    END
  END axi_master_aw_prot[0]
  PIN axi_master_aw_region[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 48.7125 0.5100 48.7875 ;
    END
  END axi_master_aw_region[3]
  PIN axi_master_aw_region[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 49.0125 0.5100 49.0875 ;
    END
  END axi_master_aw_region[2]
  PIN axi_master_aw_region[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 49.3125 0.5100 49.3875 ;
    END
  END axi_master_aw_region[1]
  PIN axi_master_aw_region[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 49.6125 0.5100 49.6875 ;
    END
  END axi_master_aw_region[0]
  PIN axi_master_aw_len[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 49.9125 0.5100 49.9875 ;
    END
  END axi_master_aw_len[7]
  PIN axi_master_aw_len[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 50.2125 0.5100 50.2875 ;
    END
  END axi_master_aw_len[6]
  PIN axi_master_aw_len[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 50.5125 0.5100 50.5875 ;
    END
  END axi_master_aw_len[5]
  PIN axi_master_aw_len[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 50.8125 0.5100 50.8875 ;
    END
  END axi_master_aw_len[4]
  PIN axi_master_aw_len[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 51.1125 0.5100 51.1875 ;
    END
  END axi_master_aw_len[3]
  PIN axi_master_aw_len[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 51.4125 0.5100 51.4875 ;
    END
  END axi_master_aw_len[2]
  PIN axi_master_aw_len[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 51.7125 0.5100 51.7875 ;
    END
  END axi_master_aw_len[1]
  PIN axi_master_aw_len[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 52.0125 0.5100 52.0875 ;
    END
  END axi_master_aw_len[0]
  PIN axi_master_aw_size[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 52.3125 0.5100 52.3875 ;
    END
  END axi_master_aw_size[2]
  PIN axi_master_aw_size[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 30.1125 0.5100 30.1875 ;
    END
  END axi_master_aw_size[1]
  PIN axi_master_aw_size[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 26.8125 0.5100 26.8875 ;
    END
  END axi_master_aw_size[0]
  PIN axi_master_aw_burst[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 52.6125 0.5100 52.6875 ;
    END
  END axi_master_aw_burst[1]
  PIN axi_master_aw_burst[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 52.9125 0.5100 52.9875 ;
    END
  END axi_master_aw_burst[0]
  PIN axi_master_aw_lock
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 53.2125 0.5100 53.2875 ;
    END
  END axi_master_aw_lock
  PIN axi_master_aw_cache[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 53.5125 0.5100 53.5875 ;
    END
  END axi_master_aw_cache[3]
  PIN axi_master_aw_cache[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 53.8125 0.5100 53.8875 ;
    END
  END axi_master_aw_cache[2]
  PIN axi_master_aw_cache[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 54.1125 0.5100 54.1875 ;
    END
  END axi_master_aw_cache[1]
  PIN axi_master_aw_cache[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 54.4125 0.5100 54.4875 ;
    END
  END axi_master_aw_cache[0]
  PIN axi_master_aw_qos[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 54.7125 0.5100 54.7875 ;
    END
  END axi_master_aw_qos[3]
  PIN axi_master_aw_qos[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 55.0125 0.5100 55.0875 ;
    END
  END axi_master_aw_qos[2]
  PIN axi_master_aw_qos[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 55.3125 0.5100 55.3875 ;
    END
  END axi_master_aw_qos[1]
  PIN axi_master_aw_qos[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 55.6125 0.5100 55.6875 ;
    END
  END axi_master_aw_qos[0]
  PIN axi_master_aw_id[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 55.9125 0.5100 55.9875 ;
    END
  END axi_master_aw_id[1]
  PIN axi_master_aw_id[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 56.2125 0.5100 56.2875 ;
    END
  END axi_master_aw_id[0]
  PIN axi_master_aw_user[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 56.5125 0.5100 56.5875 ;
    END
  END axi_master_aw_user[0]
  PIN axi_master_aw_ready
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 20.8125 0.5100 20.8875 ;
    END
  END axi_master_aw_ready
  PIN axi_master_ar_valid
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 21.5625 0.5100 21.6375 ;
    END
  END axi_master_ar_valid
  PIN axi_master_ar_addr[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 44.9625 0.5100 45.0375 ;
    END
  END axi_master_ar_addr[31]
  PIN axi_master_ar_addr[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 24.6375 66.7800 24.7125 67.2000 ;
    END
  END axi_master_ar_addr[30]
  PIN axi_master_ar_addr[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 30.7275 66.7800 30.8025 67.2000 ;
    END
  END axi_master_ar_addr[29]
  PIN axi_master_ar_addr[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 32.1975 66.7800 32.2725 67.2000 ;
    END
  END axi_master_ar_addr[28]
  PIN axi_master_ar_addr[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 32.5125 0.5100 32.5875 ;
    END
  END axi_master_ar_addr[27]
  PIN axi_master_ar_addr[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 33.4125 0.5100 33.4875 ;
    END
  END axi_master_ar_addr[26]
  PIN axi_master_ar_addr[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 32.8125 0.5100 32.8875 ;
    END
  END axi_master_ar_addr[25]
  PIN axi_master_ar_addr[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 37.6125 0.5100 37.6875 ;
    END
  END axi_master_ar_addr[24]
  PIN axi_master_ar_addr[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 39.8625 0.5100 39.9375 ;
    END
  END axi_master_ar_addr[23]
  PIN axi_master_ar_addr[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 25.6875 66.7800 25.7625 67.2000 ;
    END
  END axi_master_ar_addr[22]
  PIN axi_master_ar_addr[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 34.7175 66.7800 34.7925 67.2000 ;
    END
  END axi_master_ar_addr[21]
  PIN axi_master_ar_addr[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 31.5675 66.7800 31.6425 67.2000 ;
    END
  END axi_master_ar_addr[20]
  PIN axi_master_ar_addr[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 21.0675 66.7800 21.1425 67.2000 ;
    END
  END axi_master_ar_addr[19]
  PIN axi_master_ar_addr[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 31.9125 66.6900 31.9875 67.2000 ;
    END
  END axi_master_ar_addr[18]
  PIN axi_master_ar_addr[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17.7075 66.7800 17.7825 67.2000 ;
    END
  END axi_master_ar_addr[17]
  PIN axi_master_ar_addr[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 21.4875 66.7800 21.5625 67.2000 ;
    END
  END axi_master_ar_addr[16]
  PIN axi_master_ar_addr[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14.9775 66.7800 15.0525 67.2000 ;
    END
  END axi_master_ar_addr[15]
  PIN axi_master_ar_addr[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 20.0175 66.7800 20.0925 67.2000 ;
    END
  END axi_master_ar_addr[14]
  PIN axi_master_ar_addr[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16.8675 66.7800 16.9425 67.2000 ;
    END
  END axi_master_ar_addr[13]
  PIN axi_master_ar_addr[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 25.0575 66.7800 25.1325 67.2000 ;
    END
  END axi_master_ar_addr[12]
  PIN axi_master_ar_addr[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12.6675 66.7800 12.7425 67.2000 ;
    END
  END axi_master_ar_addr[11]
  PIN axi_master_ar_addr[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 28.4175 66.7800 28.4925 67.2000 ;
    END
  END axi_master_ar_addr[10]
  PIN axi_master_ar_addr[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 32.6175 66.7800 32.6925 67.2000 ;
    END
  END axi_master_ar_addr[9]
  PIN axi_master_ar_addr[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 34.2975 66.7800 34.3725 67.2000 ;
    END
  END axi_master_ar_addr[8]
  PIN axi_master_ar_addr[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14.5575 66.7800 14.6325 67.2000 ;
    END
  END axi_master_ar_addr[7]
  PIN axi_master_ar_addr[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 27.7875 66.7800 27.8625 67.2000 ;
    END
  END axi_master_ar_addr[6]
  PIN axi_master_ar_addr[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 19.3875 66.7800 19.4625 67.2000 ;
    END
  END axi_master_ar_addr[5]
  PIN axi_master_ar_addr[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 31.1475 66.7800 31.2225 67.2000 ;
    END
  END axi_master_ar_addr[4]
  PIN axi_master_ar_addr[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 21.9075 66.7800 21.9825 67.2000 ;
    END
  END axi_master_ar_addr[3]
  PIN axi_master_ar_addr[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 34.6125 0.5100 34.6875 ;
    END
  END axi_master_ar_addr[2]
  PIN axi_master_ar_addr[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 24.2625 0.5100 24.3375 ;
    END
  END axi_master_ar_addr[1]
  PIN axi_master_ar_addr[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 26.3625 0.5100 26.4375 ;
    END
  END axi_master_ar_addr[0]
  PIN axi_master_ar_prot[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 56.8125 0.5100 56.8875 ;
    END
  END axi_master_ar_prot[2]
  PIN axi_master_ar_prot[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 57.1125 0.5100 57.1875 ;
    END
  END axi_master_ar_prot[1]
  PIN axi_master_ar_prot[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 57.4125 0.5100 57.4875 ;
    END
  END axi_master_ar_prot[0]
  PIN axi_master_ar_region[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 57.7125 0.5100 57.7875 ;
    END
  END axi_master_ar_region[3]
  PIN axi_master_ar_region[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 58.0125 0.5100 58.0875 ;
    END
  END axi_master_ar_region[2]
  PIN axi_master_ar_region[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 58.3125 0.5100 58.3875 ;
    END
  END axi_master_ar_region[1]
  PIN axi_master_ar_region[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 58.6125 0.5100 58.6875 ;
    END
  END axi_master_ar_region[0]
  PIN axi_master_ar_len[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 58.9125 0.5100 58.9875 ;
    END
  END axi_master_ar_len[7]
  PIN axi_master_ar_len[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 59.2125 0.5100 59.2875 ;
    END
  END axi_master_ar_len[6]
  PIN axi_master_ar_len[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 59.5125 0.5100 59.5875 ;
    END
  END axi_master_ar_len[5]
  PIN axi_master_ar_len[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 59.8125 0.5100 59.8875 ;
    END
  END axi_master_ar_len[4]
  PIN axi_master_ar_len[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 60.1125 0.5100 60.1875 ;
    END
  END axi_master_ar_len[3]
  PIN axi_master_ar_len[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 60.4125 0.5100 60.4875 ;
    END
  END axi_master_ar_len[2]
  PIN axi_master_ar_len[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 60.7125 0.5100 60.7875 ;
    END
  END axi_master_ar_len[1]
  PIN axi_master_ar_len[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 61.0125 0.5100 61.0875 ;
    END
  END axi_master_ar_len[0]
  PIN axi_master_ar_size[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 61.3125 0.5100 61.3875 ;
    END
  END axi_master_ar_size[2]
  PIN axi_master_ar_size[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 30.4125 0.5100 30.4875 ;
    END
  END axi_master_ar_size[1]
  PIN axi_master_ar_size[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 27.1125 0.5100 27.1875 ;
    END
  END axi_master_ar_size[0]
  PIN axi_master_ar_burst[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 61.6125 0.5100 61.6875 ;
    END
  END axi_master_ar_burst[1]
  PIN axi_master_ar_burst[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 61.9125 0.5100 61.9875 ;
    END
  END axi_master_ar_burst[0]
  PIN axi_master_ar_lock
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 62.2125 0.5100 62.2875 ;
    END
  END axi_master_ar_lock
  PIN axi_master_ar_cache[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 62.5125 0.5100 62.5875 ;
    END
  END axi_master_ar_cache[3]
  PIN axi_master_ar_cache[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 62.8125 0.5100 62.8875 ;
    END
  END axi_master_ar_cache[2]
  PIN axi_master_ar_cache[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 63.1125 0.5100 63.1875 ;
    END
  END axi_master_ar_cache[1]
  PIN axi_master_ar_cache[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 63.4125 0.5100 63.4875 ;
    END
  END axi_master_ar_cache[0]
  PIN axi_master_ar_qos[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 63.7125 0.5100 63.7875 ;
    END
  END axi_master_ar_qos[3]
  PIN axi_master_ar_qos[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 64.0125 0.5100 64.0875 ;
    END
  END axi_master_ar_qos[2]
  PIN axi_master_ar_qos[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 64.3125 0.5100 64.3875 ;
    END
  END axi_master_ar_qos[1]
  PIN axi_master_ar_qos[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 64.6125 0.5100 64.6875 ;
    END
  END axi_master_ar_qos[0]
  PIN axi_master_ar_id[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 64.9125 0.5100 64.9875 ;
    END
  END axi_master_ar_id[1]
  PIN axi_master_ar_id[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 65.2125 0.5100 65.2875 ;
    END
  END axi_master_ar_id[0]
  PIN axi_master_ar_user[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 65.5125 0.5100 65.5875 ;
    END
  END axi_master_ar_user[0]
  PIN axi_master_ar_ready
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 23.0625 0.5100 23.1375 ;
    END
  END axi_master_ar_ready
  PIN axi_master_w_valid
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 23.0625 0.5100 23.1375 ;
    END
  END axi_master_w_valid
  PIN axi_master_w_data[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 68.3700 27.2625 68.8800 27.3375 ;
    END
  END axi_master_w_data[31]
  PIN axi_master_w_data[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 34.0125 0.0000 34.0875 0.5100 ;
    END
  END axi_master_w_data[30]
  PIN axi_master_w_data[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 31.5675 0.0000 31.6425 0.4200 ;
    END
  END axi_master_w_data[29]
  PIN axi_master_w_data[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 68.3700 26.2125 68.8800 26.2875 ;
    END
  END axi_master_w_data[28]
  PIN axi_master_w_data[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 29.8875 0.0000 29.9625 0.4200 ;
    END
  END axi_master_w_data[27]
  PIN axi_master_w_data[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 33.6675 0.0000 33.7425 0.4200 ;
    END
  END axi_master_w_data[26]
  PIN axi_master_w_data[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 68.3700 29.2125 68.8800 29.2875 ;
    END
  END axi_master_w_data[25]
  PIN axi_master_w_data[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 68.3700 28.6125 68.8800 28.6875 ;
    END
  END axi_master_w_data[24]
  PIN axi_master_w_data[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 68.3700 31.3125 68.8800 31.3875 ;
    END
  END axi_master_w_data[23]
  PIN axi_master_w_data[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 68.3700 33.1125 68.8800 33.1875 ;
    END
  END axi_master_w_data[22]
  PIN axi_master_w_data[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 68.3700 36.5625 68.8800 36.6375 ;
    END
  END axi_master_w_data[21]
  PIN axi_master_w_data[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 68.3700 34.9125 68.8800 34.9875 ;
    END
  END axi_master_w_data[20]
  PIN axi_master_w_data[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 68.3700 33.5625 68.8800 33.6375 ;
    END
  END axi_master_w_data[19]
  PIN axi_master_w_data[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 68.3700 33.4125 68.8800 33.4875 ;
    END
  END axi_master_w_data[18]
  PIN axi_master_w_data[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 38.2875 66.7800 38.3625 67.2000 ;
    END
  END axi_master_w_data[17]
  PIN axi_master_w_data[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 68.3700 35.6625 68.8800 35.7375 ;
    END
  END axi_master_w_data[16]
  PIN axi_master_w_data[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 68.3700 39.8625 68.8800 39.9375 ;
    END
  END axi_master_w_data[15]
  PIN axi_master_w_data[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 34.7625 66.6900 34.8375 67.2000 ;
    END
  END axi_master_w_data[14]
  PIN axi_master_w_data[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 35.3475 66.7800 35.4225 67.2000 ;
    END
  END axi_master_w_data[13]
  PIN axi_master_w_data[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 45.6375 66.7800 45.7125 67.2000 ;
    END
  END axi_master_w_data[12]
  PIN axi_master_w_data[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 48.3675 66.7800 48.4425 67.2000 ;
    END
  END axi_master_w_data[11]
  PIN axi_master_w_data[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 45.5625 66.6900 45.6375 67.2000 ;
    END
  END axi_master_w_data[10]
  PIN axi_master_w_data[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 37.6575 66.7800 37.7325 67.2000 ;
    END
  END axi_master_w_data[9]
  PIN axi_master_w_data[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 48.4125 66.6900 48.4875 67.2000 ;
    END
  END axi_master_w_data[8]
  PIN axi_master_w_data[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 68.3700 32.5125 68.8800 32.5875 ;
    END
  END axi_master_w_data[7]
  PIN axi_master_w_data[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 36.6075 66.7800 36.6825 67.2000 ;
    END
  END axi_master_w_data[6]
  PIN axi_master_w_data[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 42.0675 66.7800 42.1425 67.2000 ;
    END
  END axi_master_w_data[5]
  PIN axi_master_w_data[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 68.3700 45.1125 68.8800 45.1875 ;
    END
  END axi_master_w_data[4]
  PIN axi_master_w_data[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 68.3700 43.0125 68.8800 43.0875 ;
    END
  END axi_master_w_data[3]
  PIN axi_master_w_data[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 40.8075 66.7800 40.8825 67.2000 ;
    END
  END axi_master_w_data[2]
  PIN axi_master_w_data[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 36.5625 66.6900 36.6375 67.2000 ;
    END
  END axi_master_w_data[1]
  PIN axi_master_w_data[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 68.3700 46.1625 68.8800 46.2375 ;
    END
  END axi_master_w_data[0]
  PIN axi_master_w_strb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 27.4125 0.5100 27.4875 ;
    END
  END axi_master_w_strb[3]
  PIN axi_master_w_strb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 25.7625 0.5100 25.8375 ;
    END
  END axi_master_w_strb[2]
  PIN axi_master_w_strb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 27.8625 0.5100 27.9375 ;
    END
  END axi_master_w_strb[1]
  PIN axi_master_w_strb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 28.3125 0.5100 28.3875 ;
    END
  END axi_master_w_strb[0]
  PIN axi_master_w_user[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 65.8125 0.5100 65.8875 ;
    END
  END axi_master_w_user[0]
  PIN axi_master_w_last
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 65.3625 0.5100 65.4375 ;
    END
  END axi_master_w_last
  PIN axi_master_w_ready
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 22.7625 0.5100 22.8375 ;
    END
  END axi_master_w_ready
  PIN axi_master_r_valid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 24.5625 0.5100 24.6375 ;
    END
  END axi_master_r_valid
  PIN axi_master_r_data[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 47.8125 0.5100 47.8875 ;
    END
  END axi_master_r_data[31]
  PIN axi_master_r_data[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 47.2125 0.5100 47.2875 ;
    END
  END axi_master_r_data[30]
  PIN axi_master_r_data[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 46.9125 0.5100 46.9875 ;
    END
  END axi_master_r_data[29]
  PIN axi_master_r_data[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 47.5125 0.5100 47.5875 ;
    END
  END axi_master_r_data[28]
  PIN axi_master_r_data[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 38.5125 0.5100 38.5875 ;
    END
  END axi_master_r_data[27]
  PIN axi_master_r_data[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 33.2625 0.5100 33.3375 ;
    END
  END axi_master_r_data[26]
  PIN axi_master_r_data[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 35.9625 0.5100 36.0375 ;
    END
  END axi_master_r_data[25]
  PIN axi_master_r_data[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 47.2125 0.5100 47.2875 ;
    END
  END axi_master_r_data[24]
  PIN axi_master_r_data[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 46.6125 0.5100 46.6875 ;
    END
  END axi_master_r_data[23]
  PIN axi_master_r_data[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 46.9125 0.5100 46.9875 ;
    END
  END axi_master_r_data[22]
  PIN axi_master_r_data[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 48.1125 0.5100 48.1875 ;
    END
  END axi_master_r_data[21]
  PIN axi_master_r_data[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 46.3125 0.5100 46.3875 ;
    END
  END axi_master_r_data[20]
  PIN axi_master_r_data[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 37.9125 0.5100 37.9875 ;
    END
  END axi_master_r_data[19]
  PIN axi_master_r_data[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 32.5125 0.5100 32.5875 ;
    END
  END axi_master_r_data[18]
  PIN axi_master_r_data[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 34.0125 0.5100 34.0875 ;
    END
  END axi_master_r_data[17]
  PIN axi_master_r_data[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 45.2625 0.5100 45.3375 ;
    END
  END axi_master_r_data[16]
  PIN axi_master_r_data[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 46.6125 0.5100 46.6875 ;
    END
  END axi_master_r_data[15]
  PIN axi_master_r_data[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 0.0000 46.5000 2.1225 47.1000 ;
    END
  END axi_master_r_data[14]
  PIN axi_master_r_data[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 46.1625 0.5100 46.2375 ;
    END
  END axi_master_r_data[13]
  PIN axi_master_r_data[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 46.0125 0.5100 46.0875 ;
    END
  END axi_master_r_data[12]
  PIN axi_master_r_data[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 37.1625 0.5100 37.2375 ;
    END
  END axi_master_r_data[11]
  PIN axi_master_r_data[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 31.9125 0.5100 31.9875 ;
    END
  END axi_master_r_data[10]
  PIN axi_master_r_data[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 33.5625 0.5100 33.6375 ;
    END
  END axi_master_r_data[9]
  PIN axi_master_r_data[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 44.5125 0.5100 44.5875 ;
    END
  END axi_master_r_data[8]
  PIN axi_master_r_data[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 45.8625 0.5100 45.9375 ;
    END
  END axi_master_r_data[7]
  PIN axi_master_r_data[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 45.7125 0.5100 45.7875 ;
    END
  END axi_master_r_data[6]
  PIN axi_master_r_data[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 45.5625 0.5100 45.6375 ;
    END
  END axi_master_r_data[5]
  PIN axi_master_r_data[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 44.8125 0.5100 44.8875 ;
    END
  END axi_master_r_data[4]
  PIN axi_master_r_data[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 36.2625 0.5100 36.3375 ;
    END
  END axi_master_r_data[3]
  PIN axi_master_r_data[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 30.8625 0.5100 30.9375 ;
    END
  END axi_master_r_data[2]
  PIN axi_master_r_data[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 32.0625 0.5100 32.1375 ;
    END
  END axi_master_r_data[1]
  PIN axi_master_r_data[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 43.4625 0.5100 43.5375 ;
    END
  END axi_master_r_data[0]
  PIN axi_master_r_resp[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 18.5625 0.5100 18.6375 ;
    END
  END axi_master_r_resp[1]
  PIN axi_master_r_resp[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 18.4125 0.5100 18.4875 ;
    END
  END axi_master_r_resp[0]
  PIN axi_master_r_last
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 33.8775 66.7800 33.9525 67.2000 ;
    END
  END axi_master_r_last
  PIN axi_master_r_id[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 34.4625 0.0000 34.5375 0.5100 ;
    END
  END axi_master_r_id[1]
  PIN axi_master_r_id[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 34.1625 66.6900 34.2375 67.2000 ;
    END
  END axi_master_r_id[0]
  PIN axi_master_r_user[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 34.0875 0.0000 34.1625 0.4200 ;
    END
  END axi_master_r_user[0]
  PIN axi_master_r_ready
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 23.5125 0.5100 23.5875 ;
    END
  END axi_master_r_ready
  PIN axi_master_b_valid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 20.3625 0.5100 20.4375 ;
    END
  END axi_master_b_valid
  PIN axi_master_b_resp[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 19.7625 0.5100 19.8375 ;
    END
  END axi_master_b_resp[1]
  PIN axi_master_b_resp[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 19.1625 0.5100 19.2375 ;
    END
  END axi_master_b_resp[0]
  PIN axi_master_b_id[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 34.4625 66.6900 34.5375 67.2000 ;
    END
  END axi_master_b_id[1]
  PIN axi_master_b_id[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 34.5075 0.0000 34.5825 0.4200 ;
    END
  END axi_master_b_id[0]
  PIN axi_master_b_user[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 34.4625 0.0000 34.5375 0.5100 ;
    END
  END axi_master_b_user[0]
  PIN axi_master_b_ready
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 20.0625 0.5100 20.1375 ;
    END
  END axi_master_b_ready
  OBS
    LAYER M1 ;
        RECT 0.0000 0.0000 68.8800 67.2000 ;
    LAYER M2 ;
        RECT 0.0000 0.0000 68.8800 67.2000 ;
    LAYER M3 ;
        RECT 0.0000 0.0000 68.8800 67.2000 ;
    LAYER M4 ;
        RECT 0.0000 0.0000 68.8800 67.2000 ;
    LAYER M5 ;
        RECT 0.0000 0.0000 68.8800 67.2000 ;
    LAYER M6 ;
        RECT 0.0000 0.0000 68.8800 67.2000 ;
    LAYER M7 ;
        RECT 0.0000 0.0000 68.8800 67.2000 ;
    LAYER M8 ;
        RECT 0.0000 0.0000 68.8800 67.2000 ;
  END
END adv_dbg_if


VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO apb_event_unit
  CLASS BLOCK ;
    SIZE 59.4300 BY 58.8000 ;
  FOREIGN apb_event_unit 0.000000 0.000000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 34.6125 0.5100 34.6875 ;
    END
  END clk_i
  PIN HCLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 29.2575 0.0000 29.3325 0.4200 ;
    END
  END HCLK
  PIN HRESETn
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 29.3625 0.0000 29.4375 0.5100 ;
    END
  END HRESETn
  PIN PADDR[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 29.6775 58.3800 29.7525 58.8000 ;
    END
  END PADDR[11]
  PIN PADDR[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 29.6775 0.0000 29.7525 0.4200 ;
    END
  END PADDR[10]
  PIN PADDR[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 29.6625 58.2900 29.7375 58.8000 ;
    END
  END PADDR[9]
  PIN PADDR[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 29.6625 58.2900 29.7375 58.8000 ;
    END
  END PADDR[8]
  PIN PADDR[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 29.6625 0.0000 29.7375 0.5100 ;
    END
  END PADDR[7]
  PIN PADDR[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 29.6625 0.0000 29.7375 0.5100 ;
    END
  END PADDR[6]
  PIN PADDR[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 39.7575 58.3800 39.8325 58.8000 ;
    END
  END PADDR[5]
  PIN PADDR[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 31.9875 58.3800 32.0625 58.8000 ;
    END
  END PADDR[4]
  PIN PADDR[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 25.2675 58.3800 25.3425 58.8000 ;
    END
  END PADDR[3]
  PIN PADDR[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 32.3625 0.5100 32.4375 ;
    END
  END PADDR[2]
  PIN PADDR[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 29.9625 58.2900 30.0375 58.8000 ;
    END
  END PADDR[1]
  PIN PADDR[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 29.9625 58.2900 30.0375 58.8000 ;
    END
  END PADDR[0]
  PIN PWDATA[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 58.9200 10.4625 59.4300 10.5375 ;
    END
  END PWDATA[31]
  PIN PWDATA[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 58.9200 16.9125 59.4300 16.9875 ;
    END
  END PWDATA[30]
  PIN PWDATA[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 44.5875 0.0000 44.6625 0.4200 ;
    END
  END PWDATA[29]
  PIN PWDATA[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 43.9575 0.0000 44.0325 0.4200 ;
    END
  END PWDATA[28]
  PIN PWDATA[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 38.2875 0.0000 38.3625 0.4200 ;
    END
  END PWDATA[27]
  PIN PWDATA[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 28.6275 0.0000 28.7025 0.4200 ;
    END
  END PWDATA[26]
  PIN PWDATA[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 51.9375 0.0000 52.0125 0.4200 ;
    END
  END PWDATA[25]
  PIN PWDATA[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 33.2475 0.0000 33.3225 0.4200 ;
    END
  END PWDATA[24]
  PIN PWDATA[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 23.1675 0.0000 23.2425 0.4200 ;
    END
  END PWDATA[23]
  PIN PWDATA[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 19.3875 0.0000 19.4625 0.4200 ;
    END
  END PWDATA[22]
  PIN PWDATA[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 20.3625 0.5100 20.4375 ;
    END
  END PWDATA[21]
  PIN PWDATA[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 22.6125 0.5100 22.6875 ;
    END
  END PWDATA[20]
  PIN PWDATA[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14.5575 0.0000 14.6325 0.4200 ;
    END
  END PWDATA[19]
  PIN PWDATA[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 16.4625 0.5100 16.5375 ;
    END
  END PWDATA[18]
  PIN PWDATA[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 58.9200 26.8125 59.4300 26.8875 ;
    END
  END PWDATA[17]
  PIN PWDATA[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 31.5675 0.0000 31.6425 0.4200 ;
    END
  END PWDATA[16]
  PIN PWDATA[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 58.9200 26.2125 59.4300 26.2875 ;
    END
  END PWDATA[15]
  PIN PWDATA[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 58.9200 27.4125 59.4300 27.4875 ;
    END
  END PWDATA[14]
  PIN PWDATA[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 58.9200 28.3125 59.4300 28.3875 ;
    END
  END PWDATA[13]
  PIN PWDATA[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 58.9200 35.5125 59.4300 35.5875 ;
    END
  END PWDATA[12]
  PIN PWDATA[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 58.9200 48.4125 59.4300 48.4875 ;
    END
  END PWDATA[11]
  PIN PWDATA[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 58.9200 40.9125 59.4300 40.9875 ;
    END
  END PWDATA[10]
  PIN PWDATA[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 45.6375 58.3800 45.7125 58.8000 ;
    END
  END PWDATA[9]
  PIN PWDATA[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 58.9200 49.6125 59.4300 49.6875 ;
    END
  END PWDATA[8]
  PIN PWDATA[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 32.6175 58.3800 32.6925 58.8000 ;
    END
  END PWDATA[7]
  PIN PWDATA[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 40.1775 58.3800 40.2525 58.8000 ;
    END
  END PWDATA[6]
  PIN PWDATA[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 28.6275 58.3800 28.7025 58.8000 ;
    END
  END PWDATA[5]
  PIN PWDATA[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 23.1675 58.3800 23.2425 58.8000 ;
    END
  END PWDATA[4]
  PIN PWDATA[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 39.8625 0.5100 39.9375 ;
    END
  END PWDATA[3]
  PIN PWDATA[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 19.3875 58.3800 19.4625 58.8000 ;
    END
  END PWDATA[2]
  PIN PWDATA[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14.7675 58.3800 14.8425 58.8000 ;
    END
  END PWDATA[1]
  PIN PWDATA[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 33.1125 0.5100 33.1875 ;
    END
  END PWDATA[0]
  PIN PWRITE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 25.1625 58.2900 25.2375 58.8000 ;
    END
  END PWRITE
  PIN PSEL
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 32.6625 58.2900 32.7375 58.8000 ;
    END
  END PSEL
  PIN PENABLE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 33.1125 0.5100 33.1875 ;
    END
  END PENABLE
  PIN PRDATA[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 58.9200 16.0125 59.4300 16.0875 ;
    END
  END PRDATA[31]
  PIN PRDATA[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 58.9200 20.2125 59.4300 20.2875 ;
    END
  END PRDATA[30]
  PIN PRDATA[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 58.9200 19.6125 59.4300 19.6875 ;
    END
  END PRDATA[29]
  PIN PRDATA[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 43.3275 0.0000 43.4025 0.4200 ;
    END
  END PRDATA[28]
  PIN PRDATA[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 36.8175 0.0000 36.8925 0.4200 ;
    END
  END PRDATA[27]
  PIN PRDATA[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 30.9375 0.0000 31.0125 0.4200 ;
    END
  END PRDATA[26]
  PIN PRDATA[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 58.9200 18.1125 59.4300 18.1875 ;
    END
  END PRDATA[25]
  PIN PRDATA[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 32.6175 0.0000 32.6925 0.4200 ;
    END
  END PRDATA[24]
  PIN PRDATA[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 27.1575 0.0000 27.2325 0.4200 ;
    END
  END PRDATA[23]
  PIN PRDATA[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 24.2175 0.0000 24.2925 0.4200 ;
    END
  END PRDATA[22]
  PIN PRDATA[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 24.4125 0.5100 24.4875 ;
    END
  END PRDATA[21]
  PIN PRDATA[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 24.4125 0.5100 24.4875 ;
    END
  END PRDATA[20]
  PIN PRDATA[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 20.4375 0.0000 20.5125 0.4200 ;
    END
  END PRDATA[19]
  PIN PRDATA[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 22.1175 0.0000 22.1925 0.4200 ;
    END
  END PRDATA[18]
  PIN PRDATA[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 58.9200 28.6125 59.4300 28.6875 ;
    END
  END PRDATA[17]
  PIN PRDATA[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 32.1975 0.0000 32.2725 0.4200 ;
    END
  END PRDATA[16]
  PIN PRDATA[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 58.9200 26.5125 59.4300 26.5875 ;
    END
  END PRDATA[15]
  PIN PRDATA[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 58.9200 28.0125 59.4300 28.0875 ;
    END
  END PRDATA[14]
  PIN PRDATA[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 58.9200 28.0125 59.4300 28.0875 ;
    END
  END PRDATA[13]
  PIN PRDATA[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 58.9200 36.4125 59.4300 36.4875 ;
    END
  END PRDATA[12]
  PIN PRDATA[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 58.9200 41.2125 59.4300 41.2875 ;
    END
  END PRDATA[11]
  PIN PRDATA[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 58.9200 36.4125 59.4300 36.4875 ;
    END
  END PRDATA[10]
  PIN PRDATA[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 41.0175 58.3800 41.0925 58.8000 ;
    END
  END PRDATA[9]
  PIN PRDATA[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 58.9200 41.2125 59.4300 41.2875 ;
    END
  END PRDATA[8]
  PIN PRDATA[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 37.0275 58.3800 37.1025 58.8000 ;
    END
  END PRDATA[7]
  PIN PRDATA[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 38.2875 58.3800 38.3625 58.8000 ;
    END
  END PRDATA[6]
  PIN PRDATA[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 26.5275 58.3800 26.6025 58.8000 ;
    END
  END PRDATA[5]
  PIN PRDATA[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 22.7475 58.3800 22.8225 58.8000 ;
    END
  END PRDATA[4]
  PIN PRDATA[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 22.3275 58.3800 22.4025 58.8000 ;
    END
  END PRDATA[3]
  PIN PRDATA[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 24.6375 58.3800 24.7125 58.8000 ;
    END
  END PRDATA[2]
  PIN PRDATA[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 21.6975 58.3800 21.7725 58.8000 ;
    END
  END PRDATA[1]
  PIN PRDATA[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 34.3125 0.5100 34.3875 ;
    END
  END PRDATA[0]
  PIN PREADY
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 57.8625 0.5100 57.9375 ;
    END
  END PREADY
  PIN PSLVERR
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 57.8625 0.5100 57.9375 ;
    END
  END PSLVERR
  PIN irq_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 58.9200 7.1625 59.4300 7.2375 ;
    END
  END irq_i[31]
  PIN irq_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 58.9200 15.5625 59.4300 15.6375 ;
    END
  END irq_i[30]
  PIN irq_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 46.8975 0.0000 46.9725 0.4200 ;
    END
  END irq_i[29]
  PIN irq_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 46.2675 0.0000 46.3425 0.4200 ;
    END
  END irq_i[28]
  PIN irq_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 37.4475 0.0000 37.5225 0.4200 ;
    END
  END irq_i[27]
  PIN irq_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 30.0975 0.0000 30.1725 0.4200 ;
    END
  END irq_i[26]
  PIN irq_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 53.4075 0.0000 53.4825 0.4200 ;
    END
  END irq_i[25]
  PIN irq_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 34.9275 0.0000 35.0025 0.4200 ;
    END
  END irq_i[24]
  PIN irq_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 25.0575 0.0000 25.1325 0.4200 ;
    END
  END irq_i[23]
  PIN irq_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 20.8575 0.0000 20.9325 0.4200 ;
    END
  END irq_i[22]
  PIN irq_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14.5125 0.0000 14.5875 0.5100 ;
    END
  END irq_i[21]
  PIN irq_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 21.8625 0.5100 21.9375 ;
    END
  END irq_i[20]
  PIN irq_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14.1375 0.0000 14.2125 0.4200 ;
    END
  END irq_i[19]
  PIN irq_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 15.5625 0.5100 15.6375 ;
    END
  END irq_i[18]
  PIN irq_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 36.1875 0.0000 36.2625 0.4200 ;
    END
  END irq_i[17]
  PIN irq_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 33.6675 0.0000 33.7425 0.4200 ;
    END
  END irq_i[16]
  PIN irq_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 58.9200 22.1625 59.4300 22.2375 ;
    END
  END irq_i[15]
  PIN irq_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 58.9200 21.8625 59.4300 21.9375 ;
    END
  END irq_i[14]
  PIN irq_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 58.9200 25.9125 59.4300 25.9875 ;
    END
  END irq_i[13]
  PIN irq_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 58.9200 34.4625 59.4300 34.5375 ;
    END
  END irq_i[12]
  PIN irq_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 58.9200 45.2625 59.4300 45.3375 ;
    END
  END irq_i[11]
  PIN irq_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 58.9200 38.9625 59.4300 39.0375 ;
    END
  END irq_i[10]
  PIN irq_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 46.4775 58.3800 46.5525 58.8000 ;
    END
  END irq_i[9]
  PIN irq_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 58.9200 47.3625 59.4300 47.4375 ;
    END
  END irq_i[8]
  PIN irq_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 33.4575 58.3800 33.5325 58.8000 ;
    END
  END irq_i[7]
  PIN irq_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 41.8575 58.3800 41.9325 58.8000 ;
    END
  END irq_i[6]
  PIN irq_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 30.7125 58.2900 30.7875 58.8000 ;
    END
  END irq_i[5]
  PIN irq_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 21.2775 58.3800 21.3525 58.8000 ;
    END
  END irq_i[4]
  PIN irq_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 36.8625 0.5100 36.9375 ;
    END
  END irq_i[3]
  PIN irq_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18.9675 58.3800 19.0425 58.8000 ;
    END
  END irq_i[2]
  PIN irq_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14.1375 58.3800 14.2125 58.8000 ;
    END
  END irq_i[1]
  PIN irq_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 32.6625 0.5100 32.7375 ;
    END
  END irq_i[0]
  PIN event_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 58.9200 11.3625 59.4300 11.4375 ;
    END
  END event_i[31]
  PIN event_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 58.9200 17.8125 59.4300 17.8875 ;
    END
  END event_i[30]
  PIN event_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 40.3875 0.0000 40.4625 0.4200 ;
    END
  END event_i[29]
  PIN event_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 43.4625 0.0000 43.5375 0.5100 ;
    END
  END event_i[28]
  PIN event_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 38.7075 0.0000 38.7825 0.4200 ;
    END
  END event_i[27]
  PIN event_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 31.1625 0.0000 31.2375 0.5100 ;
    END
  END event_i[26]
  PIN event_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 50.8875 0.0000 50.9625 0.4200 ;
    END
  END event_i[25]
  PIN event_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 34.5075 0.0000 34.5825 0.4200 ;
    END
  END event_i[24]
  PIN event_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 26.3175 0.0000 26.3925 0.4200 ;
    END
  END event_i[23]
  PIN event_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 19.8075 0.0000 19.8825 0.4200 ;
    END
  END event_i[22]
  PIN event_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 26.3625 0.5100 26.4375 ;
    END
  END event_i[21]
  PIN event_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 23.9625 0.5100 24.0375 ;
    END
  END event_i[20]
  PIN event_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13.5075 0.0000 13.5825 0.4200 ;
    END
  END event_i[19]
  PIN event_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 17.9625 0.5100 18.0375 ;
    END
  END event_i[18]
  PIN event_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 58.9200 32.6625 59.4300 32.7375 ;
    END
  END event_i[17]
  PIN event_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 30.7275 58.3800 30.8025 58.8000 ;
    END
  END event_i[16]
  PIN event_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 58.9200 30.2625 59.4300 30.3375 ;
    END
  END event_i[15]
  PIN event_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 58.9200 32.3625 59.4300 32.4375 ;
    END
  END event_i[14]
  PIN event_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 58.9200 30.5625 59.4300 30.6375 ;
    END
  END event_i[13]
  PIN event_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 58.9200 36.7125 59.4300 36.7875 ;
    END
  END event_i[12]
  PIN event_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 58.9200 51.5625 59.4300 51.6375 ;
    END
  END event_i[11]
  PIN event_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 58.9200 42.8625 59.4300 42.9375 ;
    END
  END event_i[10]
  PIN event_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 45.0075 58.3800 45.0825 58.8000 ;
    END
  END event_i[9]
  PIN event_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 50.0475 58.3800 50.1225 58.8000 ;
    END
  END event_i[8]
  PIN event_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 36.1875 58.3800 36.2625 58.8000 ;
    END
  END event_i[7]
  PIN event_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 38.7075 58.3800 38.7825 58.8000 ;
    END
  END event_i[6]
  PIN event_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 27.9975 58.3800 28.0725 58.8000 ;
    END
  END event_i[5]
  PIN event_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 24.8625 58.2900 24.9375 58.8000 ;
    END
  END event_i[4]
  PIN event_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 41.0625 0.5100 41.1375 ;
    END
  END event_i[3]
  PIN event_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18.3375 58.3800 18.4125 58.8000 ;
    END
  END event_i[2]
  PIN event_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15.6075 58.3800 15.6825 58.8000 ;
    END
  END event_i[1]
  PIN event_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 34.9125 0.5100 34.9875 ;
    END
  END event_i[0]
  PIN irq_o[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 14.6625 0.5100 14.7375 ;
    END
  END irq_o[31]
  PIN irq_o[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 15.1125 0.5100 15.1875 ;
    END
  END irq_o[30]
  PIN irq_o[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 14.2125 0.5100 14.2875 ;
    END
  END irq_o[29]
  PIN irq_o[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 15.5625 0.5100 15.6375 ;
    END
  END irq_o[28]
  PIN irq_o[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 16.7625 0.5100 16.8375 ;
    END
  END irq_o[27]
  PIN irq_o[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 15.2625 0.5100 15.3375 ;
    END
  END irq_o[26]
  PIN irq_o[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 15.8625 0.5100 15.9375 ;
    END
  END irq_o[25]
  PIN irq_o[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 17.0625 0.5100 17.1375 ;
    END
  END irq_o[24]
  PIN irq_o[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 19.9125 0.5100 19.9875 ;
    END
  END irq_o[23]
  PIN irq_o[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 20.6625 0.5100 20.7375 ;
    END
  END irq_o[22]
  PIN irq_o[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 19.7625 0.5100 19.8375 ;
    END
  END irq_o[21]
  PIN irq_o[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 18.7125 0.5100 18.7875 ;
    END
  END irq_o[20]
  PIN irq_o[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 12.7125 0.5100 12.7875 ;
    END
  END irq_o[19]
  PIN irq_o[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 13.0125 0.5100 13.0875 ;
    END
  END irq_o[18]
  PIN irq_o[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 13.6125 0.5100 13.6875 ;
    END
  END irq_o[17]
  PIN irq_o[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 11.8125 0.5100 11.8875 ;
    END
  END irq_o[16]
  PIN irq_o[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 26.0625 0.5100 26.1375 ;
    END
  END irq_o[15]
  PIN irq_o[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 26.6625 0.5100 26.7375 ;
    END
  END irq_o[14]
  PIN irq_o[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 27.5625 0.5100 27.6375 ;
    END
  END irq_o[13]
  PIN irq_o[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 25.1625 0.5100 25.2375 ;
    END
  END irq_o[12]
  PIN irq_o[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 22.9125 0.5100 22.9875 ;
    END
  END irq_o[11]
  PIN irq_o[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 25.4625 0.5100 25.5375 ;
    END
  END irq_o[10]
  PIN irq_o[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 24.1125 0.5100 24.1875 ;
    END
  END irq_o[9]
  PIN irq_o[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 23.3625 0.5100 23.4375 ;
    END
  END irq_o[8]
  PIN irq_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 26.3625 0.5100 26.4375 ;
    END
  END irq_o[7]
  PIN irq_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 23.6625 0.5100 23.7375 ;
    END
  END irq_o[6]
  PIN irq_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 25.4625 0.5100 25.5375 ;
    END
  END irq_o[5]
  PIN irq_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 24.7125 0.5100 24.7875 ;
    END
  END irq_o[4]
  PIN irq_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 30.5625 0.5100 30.6375 ;
    END
  END irq_o[3]
  PIN irq_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 30.8625 0.5100 30.9375 ;
    END
  END irq_o[2]
  PIN irq_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 29.3625 0.5100 29.4375 ;
    END
  END irq_o[1]
  PIN irq_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 28.3125 0.5100 28.3875 ;
    END
  END irq_o[0]
  PIN fetch_enable_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 34.0125 0.5100 34.0875 ;
    END
  END fetch_enable_i
  PIN fetch_enable_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 36.5625 0.5100 36.6375 ;
    END
  END fetch_enable_o
  PIN clk_gate_core_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 33.4125 0.5100 33.4875 ;
    END
  END clk_gate_core_o
  PIN core_busy_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 32.8125 0.5100 32.8875 ;
    END
  END core_busy_i
  OBS
    LAYER M1 ;
        RECT 0.0000 0.0000 59.4300 58.8000 ;
    LAYER M2 ;
        RECT 0.0000 0.0000 59.4300 58.8000 ;
    LAYER M3 ;
        RECT 0.0000 0.0000 59.4300 58.8000 ;
    LAYER M4 ;
        RECT 0.0000 0.0000 59.4300 58.8000 ;
    LAYER M5 ;
        RECT 0.0000 0.0000 59.4300 58.8000 ;
    LAYER M6 ;
        RECT 0.0000 0.0000 59.4300 58.8000 ;
    LAYER M7 ;
        RECT 0.0000 0.0000 59.4300 58.8000 ;
    LAYER M8 ;
        RECT 0.0000 0.0000 59.4300 58.8000 ;
  END
END apb_event_unit


VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO apb_fll_if
  CLASS BLOCK ;
    SIZE 15.5400 BY 14.7000 ;
  FOREIGN apb_fll_if 0.000000 0.000000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN HCLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 10.0125 0.5100 10.0875 ;
    END
  END HCLK
  PIN HRESETn
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 9.7125 0.5100 9.7875 ;
    END
  END HRESETn
  PIN PADDR[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7.8375 14.2800 7.9125 14.7000 ;
    END
  END PADDR[11]
  PIN PADDR[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7.7625 14.1900 7.8375 14.7000 ;
    END
  END PADDR[10]
  PIN PADDR[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 7.7625 14.1900 7.8375 14.7000 ;
    END
  END PADDR[9]
  PIN PADDR[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7.8375 0.0000 7.9125 0.4200 ;
    END
  END PADDR[8]
  PIN PADDR[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7.7625 0.0000 7.8375 0.5100 ;
    END
  END PADDR[7]
  PIN PADDR[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 7.7625 0.0000 7.8375 0.5100 ;
    END
  END PADDR[6]
  PIN PADDR[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8.6775 0.0000 8.7525 0.4200 ;
    END
  END PADDR[5]
  PIN PADDR[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6.1575 0.0000 6.2325 0.4200 ;
    END
  END PADDR[4]
  PIN PADDR[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9.7275 0.0000 9.8025 0.4200 ;
    END
  END PADDR[3]
  PIN PADDR[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9.5625 0.0000 9.6375 0.5100 ;
    END
  END PADDR[2]
  PIN PADDR[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7.4175 14.2800 7.4925 14.7000 ;
    END
  END PADDR[1]
  PIN PADDR[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7.4625 14.1900 7.5375 14.7000 ;
    END
  END PADDR[0]
  PIN PWDATA[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 3.4125 0.5100 3.4875 ;
    END
  END PWDATA[31]
  PIN PWDATA[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5.3175 0.0000 5.3925 0.4200 ;
    END
  END PWDATA[30]
  PIN PWDATA[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 15.0300 2.0625 15.5400 2.1375 ;
    END
  END PWDATA[29]
  PIN PWDATA[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13.7175 0.0000 13.7925 0.4200 ;
    END
  END PWDATA[28]
  PIN PWDATA[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 15.0300 7.0125 15.5400 7.0875 ;
    END
  END PWDATA[27]
  PIN PWDATA[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9.3075 0.0000 9.3825 0.4200 ;
    END
  END PWDATA[26]
  PIN PWDATA[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4.6875 0.0000 4.7625 0.4200 ;
    END
  END PWDATA[25]
  PIN PWDATA[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 15.0300 4.9125 15.5400 4.9875 ;
    END
  END PWDATA[24]
  PIN PWDATA[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1.5375 0.0000 1.6125 0.4200 ;
    END
  END PWDATA[23]
  PIN PWDATA[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 15.0300 3.4125 15.5400 3.4875 ;
    END
  END PWDATA[22]
  PIN PWDATA[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3.0075 0.0000 3.0825 0.4200 ;
    END
  END PWDATA[21]
  PIN PWDATA[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6.7875 0.0000 6.8625 0.4200 ;
    END
  END PWDATA[20]
  PIN PWDATA[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 15.0300 3.4125 15.5400 3.4875 ;
    END
  END PWDATA[19]
  PIN PWDATA[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1.4625 0.0000 1.5375 0.5100 ;
    END
  END PWDATA[18]
  PIN PWDATA[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6.5625 0.0000 6.6375 0.5100 ;
    END
  END PWDATA[17]
  PIN PWDATA[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8.8125 0.0000 8.8875 0.5100 ;
    END
  END PWDATA[16]
  PIN PWDATA[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3.1125 0.0000 3.1875 0.5100 ;
    END
  END PWDATA[15]
  PIN PWDATA[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12.4575 0.0000 12.5325 0.4200 ;
    END
  END PWDATA[14]
  PIN PWDATA[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5.3625 0.0000 5.4375 0.5100 ;
    END
  END PWDATA[13]
  PIN PWDATA[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 2.0625 0.5100 2.1375 ;
    END
  END PWDATA[12]
  PIN PWDATA[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10.9875 0.0000 11.0625 0.4200 ;
    END
  END PWDATA[11]
  PIN PWDATA[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 9.5625 0.0000 9.6375 0.5100 ;
    END
  END PWDATA[10]
  PIN PWDATA[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 15.0300 4.1625 15.5400 4.2375 ;
    END
  END PWDATA[9]
  PIN PWDATA[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 5.3625 0.0000 5.4375 0.5100 ;
    END
  END PWDATA[8]
  PIN PWDATA[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8.2575 0.0000 8.3325 0.4200 ;
    END
  END PWDATA[7]
  PIN PWDATA[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 15.0300 4.9125 15.5400 4.9875 ;
    END
  END PWDATA[6]
  PIN PWDATA[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 6.5625 0.0000 6.6375 0.5100 ;
    END
  END PWDATA[5]
  PIN PWDATA[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 15.0300 2.8125 15.5400 2.8875 ;
    END
  END PWDATA[4]
  PIN PWDATA[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 15.0300 1.0125 15.5400 1.0875 ;
    END
  END PWDATA[3]
  PIN PWDATA[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 15.0300 6.2625 15.5400 6.3375 ;
    END
  END PWDATA[2]
  PIN PWDATA[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10.3575 0.0000 10.4325 0.4200 ;
    END
  END PWDATA[1]
  PIN PWDATA[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 3.1125 0.5100 3.1875 ;
    END
  END PWDATA[0]
  PIN PWRITE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7.4625 0.0000 7.5375 0.5100 ;
    END
  END PWRITE
  PIN PSEL
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 7.4625 0.0000 7.5375 0.5100 ;
    END
  END PSEL
  PIN PENABLE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11.4075 0.0000 11.4825 0.4200 ;
    END
  END PENABLE
  PIN PRDATA[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 15.0300 11.3625 15.5400 11.4375 ;
    END
  END PRDATA[31]
  PIN PRDATA[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 15.0300 7.4625 15.5400 7.5375 ;
    END
  END PRDATA[30]
  PIN PRDATA[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 15.0300 7.4625 15.5400 7.5375 ;
    END
  END PRDATA[29]
  PIN PRDATA[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 15.0300 9.2625 15.5400 9.3375 ;
    END
  END PRDATA[28]
  PIN PRDATA[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9.5175 14.2800 9.5925 14.7000 ;
    END
  END PRDATA[27]
  PIN PRDATA[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12.6675 14.2800 12.7425 14.7000 ;
    END
  END PRDATA[26]
  PIN PRDATA[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8.6775 14.2800 8.7525 14.7000 ;
    END
  END PRDATA[25]
  PIN PRDATA[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8.2575 14.2800 8.3325 14.7000 ;
    END
  END PRDATA[24]
  PIN PRDATA[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13.7175 14.2800 13.7925 14.7000 ;
    END
  END PRDATA[23]
  PIN PRDATA[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9.7125 14.1900 9.7875 14.7000 ;
    END
  END PRDATA[22]
  PIN PRDATA[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 9.7125 14.1900 9.7875 14.7000 ;
    END
  END PRDATA[21]
  PIN PRDATA[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 15.0300 9.2625 15.5400 9.3375 ;
    END
  END PRDATA[20]
  PIN PRDATA[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14.1375 14.2800 14.2125 14.7000 ;
    END
  END PRDATA[19]
  PIN PRDATA[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 15.0300 9.5625 15.5400 9.6375 ;
    END
  END PRDATA[18]
  PIN PRDATA[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 15.0300 11.6625 15.5400 11.7375 ;
    END
  END PRDATA[17]
  PIN PRDATA[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9.2625 14.1900 9.3375 14.7000 ;
    END
  END PRDATA[16]
  PIN PRDATA[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12.4125 14.1900 12.4875 14.7000 ;
    END
  END PRDATA[15]
  PIN PRDATA[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 15.0300 11.3625 15.5400 11.4375 ;
    END
  END PRDATA[14]
  PIN PRDATA[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12.2475 14.2800 12.3225 14.7000 ;
    END
  END PRDATA[13]
  PIN PRDATA[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9.9375 14.2800 10.0125 14.7000 ;
    END
  END PRDATA[12]
  PIN PRDATA[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 12.2625 14.1900 12.3375 14.7000 ;
    END
  END PRDATA[11]
  PIN PRDATA[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 15.0300 7.1625 15.5400 7.2375 ;
    END
  END PRDATA[10]
  PIN PRDATA[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 15.0300 8.9625 15.5400 9.0375 ;
    END
  END PRDATA[9]
  PIN PRDATA[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 15.0300 9.5625 15.5400 9.6375 ;
    END
  END PRDATA[8]
  PIN PRDATA[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 15.0300 5.3625 15.5400 5.4375 ;
    END
  END PRDATA[7]
  PIN PRDATA[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10.1625 14.1900 10.2375 14.7000 ;
    END
  END PRDATA[6]
  PIN PRDATA[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 15.0300 7.7625 15.5400 7.8375 ;
    END
  END PRDATA[5]
  PIN PRDATA[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8.2125 14.1900 8.2875 14.7000 ;
    END
  END PRDATA[4]
  PIN PRDATA[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 15.0300 9.8625 15.5400 9.9375 ;
    END
  END PRDATA[3]
  PIN PRDATA[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 8.2125 14.1900 8.2875 14.7000 ;
    END
  END PRDATA[2]
  PIN PRDATA[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8.5125 14.1900 8.5875 14.7000 ;
    END
  END PRDATA[1]
  PIN PRDATA[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8.8125 14.1900 8.8875 14.7000 ;
    END
  END PRDATA[0]
  PIN PREADY
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 6.8625 0.5100 6.9375 ;
    END
  END PREADY
  PIN PSLVERR
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 15.0300 1.3125 15.5400 1.3875 ;
    END
  END PSLVERR
  PIN fll1_req
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 5.5125 0.5100 5.5875 ;
    END
  END fll1_req
  PIN fll1_wrn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 11.3625 0.0000 11.4375 0.5100 ;
    END
  END fll1_wrn
  PIN fll1_add[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10.6125 0.0000 10.6875 0.5100 ;
    END
  END fll1_add[1]
  PIN fll1_add[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9.2625 0.0000 9.3375 0.5100 ;
    END
  END fll1_add[0]
  PIN fll1_data[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 3.4125 0.5100 3.4875 ;
    END
  END fll1_data[31]
  PIN fll1_data[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5.9625 0.0000 6.0375 0.5100 ;
    END
  END fll1_data[30]
  PIN fll1_data[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13.7625 0.0000 13.8375 0.5100 ;
    END
  END fll1_data[29]
  PIN fll1_data[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13.0875 0.0000 13.1625 0.4200 ;
    END
  END fll1_data[28]
  PIN fll1_data[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 15.0300 6.8625 15.5400 6.9375 ;
    END
  END fll1_data[27]
  PIN fll1_data[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 9.1125 0.0000 9.1875 0.5100 ;
    END
  END fll1_data[26]
  PIN fll1_data[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5.0625 0.0000 5.1375 0.5100 ;
    END
  END fll1_data[25]
  PIN fll1_data[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 15.0300 4.6125 15.5400 4.6875 ;
    END
  END fll1_data[24]
  PIN fll1_data[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2.3775 0.0000 2.4525 0.4200 ;
    END
  END fll1_data[23]
  PIN fll1_data[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 15.0300 3.1125 15.5400 3.1875 ;
    END
  END fll1_data[22]
  PIN fll1_data[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 2.8125 0.5100 2.8875 ;
    END
  END fll1_data[21]
  PIN fll1_data[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5.7375 0.0000 5.8125 0.4200 ;
    END
  END fll1_data[20]
  PIN fll1_data[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 15.0300 3.7125 15.5400 3.7875 ;
    END
  END fll1_data[19]
  PIN fll1_data[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 1.3125 0.0000 1.3875 0.5100 ;
    END
  END fll1_data[18]
  PIN fll1_data[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6.8625 0.0000 6.9375 0.5100 ;
    END
  END fll1_data[17]
  PIN fll1_data[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 8.6625 0.0000 8.7375 0.5100 ;
    END
  END fll1_data[16]
  PIN fll1_data[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3.4275 0.0000 3.5025 0.4200 ;
    END
  END fll1_data[15]
  PIN fll1_data[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12.8625 0.0000 12.9375 0.5100 ;
    END
  END fll1_data[14]
  PIN fll1_data[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 5.9625 0.0000 6.0375 0.5100 ;
    END
  END fll1_data[13]
  PIN fll1_data[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 1.6125 0.0000 1.6875 0.5100 ;
    END
  END fll1_data[12]
  PIN fll1_data[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 10.7625 0.0000 10.8375 0.5100 ;
    END
  END fll1_data[11]
  PIN fll1_data[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10.1625 0.0000 10.2375 0.5100 ;
    END
  END fll1_data[10]
  PIN fll1_data[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11.8275 0.0000 11.9025 0.4200 ;
    END
  END fll1_data[9]
  PIN fll1_data[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 5.0625 0.0000 5.1375 0.5100 ;
    END
  END fll1_data[8]
  PIN fll1_data[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8.2125 0.0000 8.2875 0.5100 ;
    END
  END fll1_data[7]
  PIN fll1_data[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 15.0300 4.6125 15.5400 4.6875 ;
    END
  END fll1_data[6]
  PIN fll1_data[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 6.8625 0.0000 6.9375 0.5100 ;
    END
  END fll1_data[5]
  PIN fll1_data[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 15.0300 2.8125 15.5400 2.8875 ;
    END
  END fll1_data[4]
  PIN fll1_data[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 15.0300 1.3125 15.5400 1.3875 ;
    END
  END fll1_data[3]
  PIN fll1_data[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 15.0300 5.5125 15.5400 5.5875 ;
    END
  END fll1_data[2]
  PIN fll1_data[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10.9125 0.0000 10.9875 0.5100 ;
    END
  END fll1_data[1]
  PIN fll1_data[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 3.7125 0.5100 3.7875 ;
    END
  END fll1_data[0]
  PIN fll1_ack
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 10.3125 0.5100 10.3875 ;
    END
  END fll1_ack
  PIN fll1_r_data[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 15.0300 11.0625 15.5400 11.1375 ;
    END
  END fll1_r_data[31]
  PIN fll1_r_data[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 15.0300 7.7625 15.5400 7.8375 ;
    END
  END fll1_r_data[30]
  PIN fll1_r_data[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 15.0300 8.0625 15.5400 8.1375 ;
    END
  END fll1_r_data[29]
  PIN fll1_r_data[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 15.0300 8.9625 15.5400 9.0375 ;
    END
  END fll1_r_data[28]
  PIN fll1_r_data[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 8.5125 14.1900 8.5875 14.7000 ;
    END
  END fll1_r_data[27]
  PIN fll1_r_data[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13.9125 14.1900 13.9875 14.7000 ;
    END
  END fll1_r_data[26]
  PIN fll1_r_data[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 10.0125 14.1900 10.0875 14.7000 ;
    END
  END fll1_r_data[25]
  PIN fll1_r_data[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 9.4125 14.1900 9.4875 14.7000 ;
    END
  END fll1_r_data[24]
  PIN fll1_r_data[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 15.0300 13.7625 15.5400 13.8375 ;
    END
  END fll1_r_data[23]
  PIN fll1_r_data[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 15.0300 8.6625 15.5400 8.7375 ;
    END
  END fll1_r_data[22]
  PIN fll1_r_data[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10.9875 14.2800 11.0625 14.7000 ;
    END
  END fll1_r_data[21]
  PIN fll1_r_data[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 15.0300 8.6625 15.5400 8.7375 ;
    END
  END fll1_r_data[20]
  PIN fll1_r_data[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 15.0300 13.1625 15.5400 13.2375 ;
    END
  END fll1_r_data[19]
  PIN fll1_r_data[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 15.0300 9.8625 15.5400 9.9375 ;
    END
  END fll1_r_data[18]
  PIN fll1_r_data[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 15.0300 11.9625 15.5400 12.0375 ;
    END
  END fll1_r_data[17]
  PIN fll1_r_data[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10.5675 14.2800 10.6425 14.7000 ;
    END
  END fll1_r_data[16]
  PIN fll1_r_data[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11.2125 14.1900 11.2875 14.7000 ;
    END
  END fll1_r_data[15]
  PIN fll1_r_data[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 15.0300 11.0625 15.5400 11.1375 ;
    END
  END fll1_r_data[14]
  PIN fll1_r_data[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13.4625 14.1900 13.5375 14.7000 ;
    END
  END fll1_r_data[13]
  PIN fll1_r_data[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10.9125 14.1900 10.9875 14.7000 ;
    END
  END fll1_r_data[12]
  PIN fll1_r_data[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 15.0300 11.9625 15.5400 12.0375 ;
    END
  END fll1_r_data[11]
  PIN fll1_r_data[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 15.0300 8.0625 15.5400 8.1375 ;
    END
  END fll1_r_data[10]
  PIN fll1_r_data[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 15.0300 8.3625 15.5400 8.4375 ;
    END
  END fll1_r_data[9]
  PIN fll1_r_data[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 15.0300 10.1625 15.5400 10.2375 ;
    END
  END fll1_r_data[8]
  PIN fll1_r_data[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 15.0300 5.6625 15.5400 5.7375 ;
    END
  END fll1_r_data[7]
  PIN fll1_r_data[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11.4075 14.2800 11.4825 14.7000 ;
    END
  END fll1_r_data[6]
  PIN fll1_r_data[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 15.0300 8.3625 15.5400 8.4375 ;
    END
  END fll1_r_data[5]
  PIN fll1_r_data[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 13.4175 6.9000 15.5400 7.5000 ;
    END
  END fll1_r_data[4]
  PIN fll1_r_data[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 15.0300 10.1625 15.5400 10.2375 ;
    END
  END fll1_r_data[3]
  PIN fll1_r_data[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9.0975 14.2800 9.1725 14.7000 ;
    END
  END fll1_r_data[2]
  PIN fll1_r_data[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 10.3125 14.1900 10.3875 14.7000 ;
    END
  END fll1_r_data[1]
  PIN fll1_r_data[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 8.8125 14.1900 8.8875 14.7000 ;
    END
  END fll1_r_data[0]
  PIN fll1_lock
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3.8475 14.2800 3.9225 14.7000 ;
    END
  END fll1_lock
  PIN fll2_req
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 6.4125 0.5100 6.4875 ;
    END
  END fll2_req
  PIN fll2_wrn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6.2625 0.0000 6.3375 0.5100 ;
    END
  END fll2_wrn
  PIN fll2_add[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 10.3125 0.0000 10.3875 0.5100 ;
    END
  END fll2_add[1]
  PIN fll2_add[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9.8625 0.0000 9.9375 0.5100 ;
    END
  END fll2_add[0]
  PIN fll2_data[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 3.1125 0.5100 3.1875 ;
    END
  END fll2_data[31]
  PIN fll2_data[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4.7625 0.0000 4.8375 0.5100 ;
    END
  END fll2_data[30]
  PIN fll2_data[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 15.0300 2.5125 15.5400 2.5875 ;
    END
  END fll2_data[29]
  PIN fll2_data[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14.1375 0.0000 14.2125 0.4200 ;
    END
  END fll2_data[28]
  PIN fll2_data[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 15.0300 6.7125 15.5400 6.7875 ;
    END
  END fll2_data[27]
  PIN fll2_data[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 9.8625 0.0000 9.9375 0.5100 ;
    END
  END fll2_data[26]
  PIN fll2_data[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4.0575 0.0000 4.1325 0.4200 ;
    END
  END fll2_data[25]
  PIN fll2_data[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 15.0300 5.2125 15.5400 5.2875 ;
    END
  END fll2_data[24]
  PIN fll2_data[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1.3125 0.5100 1.3875 ;
    END
  END fll2_data[23]
  PIN fll2_data[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 15.0300 3.1125 15.5400 3.1875 ;
    END
  END fll2_data[22]
  PIN fll2_data[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3.4125 0.0000 3.4875 0.5100 ;
    END
  END fll2_data[21]
  PIN fll2_data[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7.4175 0.0000 7.4925 0.4200 ;
    END
  END fll2_data[20]
  PIN fll2_data[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 15.0300 3.7125 15.5400 3.7875 ;
    END
  END fll2_data[19]
  PIN fll2_data[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2.2125 0.0000 2.2875 0.5100 ;
    END
  END fll2_data[18]
  PIN fll2_data[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7.1625 0.0000 7.2375 0.5100 ;
    END
  END fll2_data[17]
  PIN fll2_data[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8.5125 0.0000 8.5875 0.5100 ;
    END
  END fll2_data[16]
  PIN fll2_data[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2.8125 0.0000 2.8875 0.5100 ;
    END
  END fll2_data[15]
  PIN fll2_data[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12.4125 0.0000 12.4875 0.5100 ;
    END
  END fll2_data[14]
  PIN fll2_data[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 4.7625 0.0000 4.8375 0.5100 ;
    END
  END fll2_data[13]
  PIN fll2_data[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 2.8125 0.5100 2.8875 ;
    END
  END fll2_data[12]
  PIN fll2_data[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 11.0625 0.0000 11.1375 0.5100 ;
    END
  END fll2_data[11]
  PIN fll2_data[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 8.3625 0.0000 8.4375 0.5100 ;
    END
  END fll2_data[10]
  PIN fll2_data[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 15.0300 4.3125 15.5400 4.3875 ;
    END
  END fll2_data[9]
  PIN fll2_data[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5.6625 0.0000 5.7375 0.5100 ;
    END
  END fll2_data[8]
  PIN fll2_data[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 8.0625 0.0000 8.1375 0.5100 ;
    END
  END fll2_data[7]
  PIN fll2_data[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 15.0300 4.0125 15.5400 4.0875 ;
    END
  END fll2_data[6]
  PIN fll2_data[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 7.1625 0.0000 7.2375 0.5100 ;
    END
  END fll2_data[5]
  PIN fll2_data[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 12.8625 0.0000 12.9375 0.5100 ;
    END
  END fll2_data[4]
  PIN fll2_data[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14.6625 0.0000 14.7375 0.5100 ;
    END
  END fll2_data[3]
  PIN fll2_data[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 15.0300 6.5625 15.5400 6.6375 ;
    END
  END fll2_data[2]
  PIN fll2_data[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11.2125 0.0000 11.2875 0.5100 ;
    END
  END fll2_data[1]
  PIN fll2_data[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 2.5125 0.5100 2.5875 ;
    END
  END fll2_data[0]
  PIN fll2_ack
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 12.1125 0.5100 12.1875 ;
    END
  END fll2_ack
  PIN fll2_r_data[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 15.0300 10.7625 15.5400 10.8375 ;
    END
  END fll2_r_data[31]
  PIN fll2_r_data[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 15.0300 6.4125 15.5400 6.4875 ;
    END
  END fll2_r_data[30]
  PIN fll2_r_data[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 15.0300 5.9625 15.5400 6.0375 ;
    END
  END fll2_r_data[29]
  PIN fll2_r_data[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 15.0300 10.4625 15.5400 10.5375 ;
    END
  END fll2_r_data[28]
  PIN fll2_r_data[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 9.1125 14.1900 9.1875 14.7000 ;
    END
  END fll2_r_data[27]
  PIN fll2_r_data[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13.0875 14.2800 13.1625 14.7000 ;
    END
  END fll2_r_data[26]
  PIN fll2_r_data[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10.4625 14.1900 10.5375 14.7000 ;
    END
  END fll2_r_data[25]
  PIN fll2_r_data[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6.9975 14.2800 7.0725 14.7000 ;
    END
  END fll2_r_data[24]
  PIN fll2_r_data[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14.2125 14.1900 14.2875 14.7000 ;
    END
  END fll2_r_data[23]
  PIN fll2_r_data[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 10.6125 14.1900 10.6875 14.7000 ;
    END
  END fll2_r_data[22]
  PIN fll2_r_data[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 10.9125 14.1900 10.9875 14.7000 ;
    END
  END fll2_r_data[21]
  PIN fll2_r_data[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 15.0300 10.4625 15.5400 10.5375 ;
    END
  END fll2_r_data[20]
  PIN fll2_r_data[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 15.0300 12.8625 15.5400 12.9375 ;
    END
  END fll2_r_data[19]
  PIN fll2_r_data[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11.8275 14.2800 11.9025 14.7000 ;
    END
  END fll2_r_data[18]
  PIN fll2_r_data[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 15.0300 12.2625 15.5400 12.3375 ;
    END
  END fll2_r_data[17]
  PIN fll2_r_data[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11.5125 14.1900 11.5875 14.7000 ;
    END
  END fll2_r_data[16]
  PIN fll2_r_data[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11.9625 14.1900 12.0375 14.7000 ;
    END
  END fll2_r_data[15]
  PIN fll2_r_data[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 15.0300 10.7625 15.5400 10.8375 ;
    END
  END fll2_r_data[14]
  PIN fll2_r_data[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12.7125 14.1900 12.7875 14.7000 ;
    END
  END fll2_r_data[13]
  PIN fll2_r_data[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 11.2125 14.1900 11.2875 14.7000 ;
    END
  END fll2_r_data[12]
  PIN fll2_r_data[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13.0125 14.1900 13.0875 14.7000 ;
    END
  END fll2_r_data[11]
  PIN fll2_r_data[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 15.0300 6.1125 15.5400 6.1875 ;
    END
  END fll2_r_data[10]
  PIN fll2_r_data[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 15.0300 11.6625 15.5400 11.7375 ;
    END
  END fll2_r_data[9]
  PIN fll2_r_data[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 15.0300 12.5625 15.5400 12.6375 ;
    END
  END fll2_r_data[8]
  PIN fll2_r_data[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 15.0300 5.8125 15.5400 5.8875 ;
    END
  END fll2_r_data[7]
  PIN fll2_r_data[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 11.5125 14.1900 11.5875 14.7000 ;
    END
  END fll2_r_data[6]
  PIN fll2_r_data[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 15.0300 12.2625 15.5400 12.3375 ;
    END
  END fll2_r_data[5]
  PIN fll2_r_data[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7.1625 14.1900 7.2375 14.7000 ;
    END
  END fll2_r_data[4]
  PIN fll2_r_data[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 13.0125 14.1900 13.0875 14.7000 ;
    END
  END fll2_r_data[3]
  PIN fll2_r_data[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 7.4625 14.1900 7.5375 14.7000 ;
    END
  END fll2_r_data[2]
  PIN fll2_r_data[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 7.1625 14.1900 7.2375 14.7000 ;
    END
  END fll2_r_data[1]
  PIN fll2_r_data[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 11.8125 14.1900 11.8875 14.7000 ;
    END
  END fll2_r_data[0]
  PIN fll2_lock
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3.8625 14.1900 3.9375 14.7000 ;
    END
  END fll2_lock
  OBS
    LAYER M1 ;
        RECT 0.0000 0.0000 15.5400 14.7000 ;
    LAYER M2 ;
        RECT 0.0000 0.0000 15.5400 14.7000 ;
    LAYER M3 ;
        RECT 0.0000 0.0000 15.5400 14.7000 ;
    LAYER M4 ;
        RECT 0.0000 0.0000 15.5400 14.7000 ;
    LAYER M5 ;
        RECT 0.0000 0.0000 15.5400 14.7000 ;
    LAYER M6 ;
        RECT 0.0000 0.0000 15.5400 14.7000 ;
    LAYER M7 ;
        RECT 0.0000 0.0000 15.5400 14.7000 ;
    LAYER M8 ;
        RECT 0.0000 0.0000 15.5400 14.7000 ;
  END
END apb_fll_if


VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO apb_i2c
  CLASS BLOCK ;
    SIZE 35.7000 BY 34.6500 ;
  FOREIGN apb_i2c 0.000000 0.000000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN HCLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 17.6625 0.5100 17.7375 ;
    END
  END HCLK
  PIN HRESETn
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17.0775 34.2300 17.1525 34.6500 ;
    END
  END HRESETn
  PIN PADDR[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17.9175 34.2300 17.9925 34.6500 ;
    END
  END PADDR[11]
  PIN PADDR[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17.8125 34.1400 17.8875 34.6500 ;
    END
  END PADDR[10]
  PIN PADDR[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 17.8125 34.1400 17.8875 34.6500 ;
    END
  END PADDR[9]
  PIN PADDR[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17.9175 0.0000 17.9925 0.4200 ;
    END
  END PADDR[8]
  PIN PADDR[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17.8125 0.0000 17.8875 0.5100 ;
    END
  END PADDR[7]
  PIN PADDR[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 17.8125 0.0000 17.8875 0.5100 ;
    END
  END PADDR[6]
  PIN PADDR[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 20.4375 0.0000 20.5125 0.4200 ;
    END
  END PADDR[5]
  PIN PADDR[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 21.6975 0.0000 21.7725 0.4200 ;
    END
  END PADDR[4]
  PIN PADDR[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 20.3625 0.0000 20.4375 0.5100 ;
    END
  END PADDR[3]
  PIN PADDR[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 22.1175 0.0000 22.1925 0.4200 ;
    END
  END PADDR[2]
  PIN PADDR[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17.4975 34.2300 17.5725 34.6500 ;
    END
  END PADDR[1]
  PIN PADDR[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17.5125 34.1400 17.5875 34.6500 ;
    END
  END PADDR[0]
  PIN PWDATA[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18.1125 34.1400 18.1875 34.6500 ;
    END
  END PWDATA[31]
  PIN PWDATA[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 17.5125 34.1400 17.5875 34.6500 ;
    END
  END PWDATA[30]
  PIN PWDATA[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 18.1125 34.1400 18.1875 34.6500 ;
    END
  END PWDATA[29]
  PIN PWDATA[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17.4975 0.0000 17.5725 0.4200 ;
    END
  END PWDATA[28]
  PIN PWDATA[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17.5125 0.0000 17.5875 0.5100 ;
    END
  END PWDATA[27]
  PIN PWDATA[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 17.5125 0.0000 17.5875 0.5100 ;
    END
  END PWDATA[26]
  PIN PWDATA[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 18.1125 0.0000 18.1875 0.5100 ;
    END
  END PWDATA[25]
  PIN PWDATA[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18.3375 34.2300 18.4125 34.6500 ;
    END
  END PWDATA[24]
  PIN PWDATA[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 17.2125 0.5100 17.2875 ;
    END
  END PWDATA[23]
  PIN PWDATA[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 17.2125 0.5100 17.2875 ;
    END
  END PWDATA[22]
  PIN PWDATA[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17.2125 34.1400 17.2875 34.6500 ;
    END
  END PWDATA[21]
  PIN PWDATA[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18.4125 34.1400 18.4875 34.6500 ;
    END
  END PWDATA[20]
  PIN PWDATA[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 17.2125 34.1400 17.2875 34.6500 ;
    END
  END PWDATA[19]
  PIN PWDATA[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 18.4125 34.1400 18.4875 34.6500 ;
    END
  END PWDATA[18]
  PIN PWDATA[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 35.1900 17.2125 35.7000 17.2875 ;
    END
  END PWDATA[17]
  PIN PWDATA[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 35.1900 17.2125 35.7000 17.2875 ;
    END
  END PWDATA[16]
  PIN PWDATA[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 23.1675 34.2300 23.2425 34.6500 ;
    END
  END PWDATA[15]
  PIN PWDATA[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 22.1175 34.2300 22.1925 34.6500 ;
    END
  END PWDATA[14]
  PIN PWDATA[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 25.2675 34.2300 25.3425 34.6500 ;
    END
  END PWDATA[13]
  PIN PWDATA[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 35.1900 26.6625 35.7000 26.7375 ;
    END
  END PWDATA[12]
  PIN PWDATA[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 35.1900 27.8625 35.7000 27.9375 ;
    END
  END PWDATA[11]
  PIN PWDATA[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 35.1900 24.5625 35.7000 24.6375 ;
    END
  END PWDATA[10]
  PIN PWDATA[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 35.1900 27.5625 35.7000 27.6375 ;
    END
  END PWDATA[9]
  PIN PWDATA[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 35.1900 22.4625 35.7000 22.5375 ;
    END
  END PWDATA[8]
  PIN PWDATA[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 35.1900 16.1625 35.7000 16.2375 ;
    END
  END PWDATA[7]
  PIN PWDATA[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 35.1900 14.0625 35.7000 14.1375 ;
    END
  END PWDATA[6]
  PIN PWDATA[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 18.7125 0.0000 18.7875 0.5100 ;
    END
  END PWDATA[5]
  PIN PWDATA[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11.4075 0.0000 11.4825 0.4200 ;
    END
  END PWDATA[4]
  PIN PWDATA[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11.3625 0.0000 11.4375 0.5100 ;
    END
  END PWDATA[3]
  PIN PWDATA[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 30.5175 0.0000 30.5925 0.4200 ;
    END
  END PWDATA[2]
  PIN PWDATA[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 29.0475 0.0000 29.1225 0.4200 ;
    END
  END PWDATA[1]
  PIN PWDATA[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 11.2125 0.0000 11.2875 0.5100 ;
    END
  END PWDATA[0]
  PIN PWRITE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 21.0675 0.0000 21.1425 0.4200 ;
    END
  END PWRITE
  PIN PSEL
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 20.6625 0.0000 20.7375 0.5100 ;
    END
  END PSEL
  PIN PENABLE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 20.8125 0.0000 20.8875 0.5100 ;
    END
  END PENABLE
  PIN PRDATA[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 4.6125 0.0000 4.6875 0.5100 ;
    END
  END PRDATA[31]
  PIN PRDATA[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 4.3125 0.0000 4.3875 0.5100 ;
    END
  END PRDATA[30]
  PIN PRDATA[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 4.0125 0.0000 4.0875 0.5100 ;
    END
  END PRDATA[29]
  PIN PRDATA[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 3.7125 0.0000 3.7875 0.5100 ;
    END
  END PRDATA[28]
  PIN PRDATA[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 3.4125 0.0000 3.4875 0.5100 ;
    END
  END PRDATA[27]
  PIN PRDATA[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 3.1125 0.0000 3.1875 0.5100 ;
    END
  END PRDATA[26]
  PIN PRDATA[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 2.8125 0.0000 2.8875 0.5100 ;
    END
  END PRDATA[25]
  PIN PRDATA[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 2.5125 0.0000 2.5875 0.5100 ;
    END
  END PRDATA[24]
  PIN PRDATA[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 2.2125 0.0000 2.2875 0.5100 ;
    END
  END PRDATA[23]
  PIN PRDATA[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 1.9125 0.0000 1.9875 0.5100 ;
    END
  END PRDATA[22]
  PIN PRDATA[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 1.6125 0.0000 1.6875 0.5100 ;
    END
  END PRDATA[21]
  PIN PRDATA[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 1.3125 0.0000 1.3875 0.5100 ;
    END
  END PRDATA[20]
  PIN PRDATA[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 1.0125 0.0000 1.0875 0.5100 ;
    END
  END PRDATA[19]
  PIN PRDATA[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1.0125 0.0000 1.0875 0.5100 ;
    END
  END PRDATA[18]
  PIN PRDATA[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1.3125 0.0000 1.3875 0.5100 ;
    END
  END PRDATA[17]
  PIN PRDATA[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1.6125 0.0000 1.6875 0.5100 ;
    END
  END PRDATA[16]
  PIN PRDATA[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 22.5375 34.2300 22.6125 34.6500 ;
    END
  END PRDATA[15]
  PIN PRDATA[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 24.0075 34.2300 24.0825 34.6500 ;
    END
  END PRDATA[14]
  PIN PRDATA[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 24.8475 34.2300 24.9225 34.6500 ;
    END
  END PRDATA[13]
  PIN PRDATA[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 26.3175 34.2300 26.3925 34.6500 ;
    END
  END PRDATA[12]
  PIN PRDATA[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 35.1900 28.1625 35.7000 28.2375 ;
    END
  END PRDATA[11]
  PIN PRDATA[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 35.1900 26.3625 35.7000 26.4375 ;
    END
  END PRDATA[10]
  PIN PRDATA[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 35.1900 28.1625 35.7000 28.2375 ;
    END
  END PRDATA[9]
  PIN PRDATA[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 35.1900 21.8625 35.7000 21.9375 ;
    END
  END PRDATA[8]
  PIN PRDATA[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 19.3875 0.0000 19.4625 0.4200 ;
    END
  END PRDATA[7]
  PIN PRDATA[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18.9675 0.0000 19.0425 0.4200 ;
    END
  END PRDATA[6]
  PIN PRDATA[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18.5475 0.0000 18.6225 0.4200 ;
    END
  END PRDATA[5]
  PIN PRDATA[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18.7125 0.0000 18.7875 0.5100 ;
    END
  END PRDATA[4]
  PIN PRDATA[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 19.8075 0.0000 19.8825 0.4200 ;
    END
  END PRDATA[3]
  PIN PRDATA[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 21.4125 0.0000 21.4875 0.5100 ;
    END
  END PRDATA[2]
  PIN PRDATA[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 21.7125 0.0000 21.7875 0.5100 ;
    END
  END PRDATA[1]
  PIN PRDATA[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18.1125 0.0000 18.1875 0.5100 ;
    END
  END PRDATA[0]
  PIN PREADY
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 34.5075 0.0000 34.5825 0.4200 ;
    END
  END PREADY
  PIN PSLVERR
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1.9125 0.0000 1.9875 0.5100 ;
    END
  END PSLVERR
  PIN interrupt_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4.8975 0.0000 4.9725 0.4200 ;
    END
  END interrupt_o
  PIN scl_pad_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 19.5975 34.2300 19.6725 34.6500 ;
    END
  END scl_pad_i
  PIN scl_pad_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2.2125 0.0000 2.2875 0.5100 ;
    END
  END scl_pad_o
  PIN scl_padoen_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16.0275 34.2300 16.1025 34.6500 ;
    END
  END scl_padoen_o
  PIN sda_pad_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9.5175 34.2300 9.5925 34.6500 ;
    END
  END sda_pad_i
  PIN sda_pad_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2.1675 0.0000 2.2425 0.4200 ;
    END
  END sda_pad_o
  PIN sda_padoen_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11.6175 34.2300 11.6925 34.6500 ;
    END
  END sda_padoen_o
  OBS
    LAYER M1 ;
        RECT 0.0000 0.0000 35.7000 34.6500 ;
    LAYER M2 ;
        RECT 0.0000 0.0000 35.7000 34.6500 ;
    LAYER M3 ;
        RECT 0.0000 0.0000 35.7000 34.6500 ;
    LAYER M4 ;
        RECT 0.0000 0.0000 35.7000 34.6500 ;
    LAYER M5 ;
        RECT 0.0000 0.0000 35.7000 34.6500 ;
    LAYER M6 ;
        RECT 0.0000 0.0000 35.7000 34.6500 ;
    LAYER M7 ;
        RECT 0.0000 0.0000 35.7000 34.6500 ;
    LAYER M8 ;
        RECT 0.0000 0.0000 35.7000 34.6500 ;
  END
END apb_i2c


VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO apb_pulpino
  CLASS BLOCK ;
    SIZE 49.3500 BY 48.3000 ;
  FOREIGN apb_pulpino 0.000000 0.000000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN HCLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 48.8400 23.6625 49.3500 23.7375 ;
    END
  END HCLK
  PIN HRESETn
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 24.8625 0.0000 24.9375 0.5100 ;
    END
  END HRESETn
  PIN PADDR[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 24.6375 47.8800 24.7125 48.3000 ;
    END
  END PADDR[11]
  PIN PADDR[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 24.6375 0.0000 24.7125 0.4200 ;
    END
  END PADDR[10]
  PIN PADDR[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 24.5625 47.7900 24.6375 48.3000 ;
    END
  END PADDR[9]
  PIN PADDR[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 24.5625 47.7900 24.6375 48.3000 ;
    END
  END PADDR[8]
  PIN PADDR[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 24.5625 0.0000 24.6375 0.5100 ;
    END
  END PADDR[7]
  PIN PADDR[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 24.5625 0.0000 24.6375 0.5100 ;
    END
  END PADDR[6]
  PIN PADDR[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15.1875 47.8800 15.2625 48.3000 ;
    END
  END PADDR[5]
  PIN PADDR[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12.8775 47.8800 12.9525 48.3000 ;
    END
  END PADDR[4]
  PIN PADDR[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16.2375 47.8800 16.3125 48.3000 ;
    END
  END PADDR[3]
  PIN PADDR[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13.7175 47.8800 13.7925 48.3000 ;
    END
  END PADDR[2]
  PIN PADDR[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 24.8625 47.7900 24.9375 48.3000 ;
    END
  END PADDR[1]
  PIN PADDR[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 24.8625 47.7900 24.9375 48.3000 ;
    END
  END PADDR[0]
  PIN PWDATA[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 27.5775 47.8800 27.6525 48.3000 ;
    END
  END PWDATA[31]
  PIN PWDATA[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 28.7625 0.5100 28.8375 ;
    END
  END PWDATA[30]
  PIN PWDATA[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 48.8400 22.4625 49.3500 22.5375 ;
    END
  END PWDATA[29]
  PIN PWDATA[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 21.5625 0.5100 21.6375 ;
    END
  END PWDATA[28]
  PIN PWDATA[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 48.8400 22.4625 49.3500 22.5375 ;
    END
  END PWDATA[27]
  PIN PWDATA[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 29.9625 0.5100 30.0375 ;
    END
  END PWDATA[26]
  PIN PWDATA[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 48.8400 27.8625 49.3500 27.9375 ;
    END
  END PWDATA[25]
  PIN PWDATA[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 48.8400 11.9625 49.3500 12.0375 ;
    END
  END PWDATA[24]
  PIN PWDATA[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 35.0625 0.5100 35.1375 ;
    END
  END PWDATA[23]
  PIN PWDATA[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 16.1625 0.5100 16.2375 ;
    END
  END PWDATA[22]
  PIN PWDATA[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 48.8400 24.5625 49.3500 24.6375 ;
    END
  END PWDATA[21]
  PIN PWDATA[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 47.1075 47.8800 47.1825 48.3000 ;
    END
  END PWDATA[20]
  PIN PWDATA[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17.4975 0.0000 17.5725 0.4200 ;
    END
  END PWDATA[19]
  PIN PWDATA[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2.3775 0.0000 2.4525 0.4200 ;
    END
  END PWDATA[18]
  PIN PWDATA[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 25.4775 0.0000 25.5525 0.4200 ;
    END
  END PWDATA[17]
  PIN PWDATA[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 41.2275 47.8800 41.3025 48.3000 ;
    END
  END PWDATA[16]
  PIN PWDATA[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 45.5625 0.5100 45.6375 ;
    END
  END PWDATA[15]
  PIN PWDATA[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 24.5625 0.5100 24.6375 ;
    END
  END PWDATA[14]
  PIN PWDATA[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 37.4625 0.0000 37.5375 0.5100 ;
    END
  END PWDATA[13]
  PIN PWDATA[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 21.2775 0.0000 21.3525 0.4200 ;
    END
  END PWDATA[12]
  PIN PWDATA[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 48.8400 14.0625 49.3500 14.1375 ;
    END
  END PWDATA[11]
  PIN PWDATA[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 48.8400 34.1625 49.3500 34.2375 ;
    END
  END PWDATA[10]
  PIN PWDATA[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16.4475 0.0000 16.5225 0.4200 ;
    END
  END PWDATA[9]
  PIN PWDATA[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 32.4075 47.8800 32.4825 48.3000 ;
    END
  END PWDATA[8]
  PIN PWDATA[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 45.5625 0.5100 45.6375 ;
    END
  END PWDATA[7]
  PIN PWDATA[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 0.0000 21.3000 2.1225 21.9000 ;
    END
  END PWDATA[6]
  PIN PWDATA[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 25.7625 0.5100 25.8375 ;
    END
  END PWDATA[5]
  PIN PWDATA[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 7.7625 0.5100 7.8375 ;
    END
  END PWDATA[4]
  PIN PWDATA[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 32.4075 0.0000 32.4825 0.4200 ;
    END
  END PWDATA[3]
  PIN PWDATA[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 25.6125 0.5100 25.6875 ;
    END
  END PWDATA[2]
  PIN PWDATA[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6.1575 47.8800 6.2325 48.3000 ;
    END
  END PWDATA[1]
  PIN PWDATA[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18.5475 47.8800 18.6225 48.3000 ;
    END
  END PWDATA[0]
  PIN PWRITE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 18.7125 47.7900 18.7875 48.3000 ;
    END
  END PWRITE
  PIN PSEL
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 19.5975 47.8800 19.6725 48.3000 ;
    END
  END PSEL
  PIN PENABLE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 19.3125 47.7900 19.3875 48.3000 ;
    END
  END PENABLE
  PIN PRDATA[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 24.0075 47.8800 24.0825 48.3000 ;
    END
  END PRDATA[31]
  PIN PRDATA[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 28.0125 0.5100 28.0875 ;
    END
  END PRDATA[30]
  PIN PRDATA[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 48.8400 20.6625 49.3500 20.7375 ;
    END
  END PRDATA[29]
  PIN PRDATA[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 17.0625 0.5100 17.1375 ;
    END
  END PRDATA[28]
  PIN PRDATA[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 31.3575 0.0000 31.4325 0.4200 ;
    END
  END PRDATA[27]
  PIN PRDATA[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 26.9625 0.5100 27.0375 ;
    END
  END PRDATA[26]
  PIN PRDATA[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 48.8400 27.5625 49.3500 27.6375 ;
    END
  END PRDATA[25]
  PIN PRDATA[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 37.6575 0.0000 37.7325 0.4200 ;
    END
  END PRDATA[24]
  PIN PRDATA[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 32.8125 0.5100 32.8875 ;
    END
  END PRDATA[23]
  PIN PRDATA[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 17.5125 0.5100 17.5875 ;
    END
  END PRDATA[22]
  PIN PRDATA[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 48.8400 26.9625 49.3500 27.0375 ;
    END
  END PRDATA[21]
  PIN PRDATA[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 37.2375 47.8800 37.3125 48.3000 ;
    END
  END PRDATA[20]
  PIN PRDATA[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 16.4625 0.5100 16.5375 ;
    END
  END PRDATA[19]
  PIN PRDATA[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 8.6625 0.5100 8.7375 ;
    END
  END PRDATA[18]
  PIN PRDATA[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 23.5875 0.0000 23.6625 0.4200 ;
    END
  END PRDATA[17]
  PIN PRDATA[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 37.8675 47.8800 37.9425 48.3000 ;
    END
  END PRDATA[16]
  PIN PRDATA[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5.1075 47.8800 5.1825 48.3000 ;
    END
  END PRDATA[15]
  PIN PRDATA[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 25.9125 0.5100 25.9875 ;
    END
  END PRDATA[14]
  PIN PRDATA[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 35.1375 0.0000 35.2125 0.4200 ;
    END
  END PRDATA[13]
  PIN PRDATA[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 23.1675 0.0000 23.2425 0.4200 ;
    END
  END PRDATA[12]
  PIN PRDATA[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 48.8400 16.4625 49.3500 16.5375 ;
    END
  END PRDATA[11]
  PIN PRDATA[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 48.8400 33.8625 49.3500 33.9375 ;
    END
  END PRDATA[10]
  PIN PRDATA[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17.0775 0.0000 17.1525 0.4200 ;
    END
  END PRDATA[9]
  PIN PRDATA[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 30.0975 47.8800 30.1725 48.3000 ;
    END
  END PRDATA[8]
  PIN PRDATA[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 43.3125 0.5100 43.3875 ;
    END
  END PRDATA[7]
  PIN PRDATA[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 21.7125 0.5100 21.7875 ;
    END
  END PRDATA[6]
  PIN PRDATA[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 20.8575 47.8800 20.9325 48.3000 ;
    END
  END PRDATA[5]
  PIN PRDATA[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 12.8625 0.5100 12.9375 ;
    END
  END PRDATA[4]
  PIN PRDATA[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 28.6275 0.0000 28.7025 0.4200 ;
    END
  END PRDATA[3]
  PIN PRDATA[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 29.0625 0.5100 29.1375 ;
    END
  END PRDATA[2]
  PIN PRDATA[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11.1975 47.8800 11.2725 48.3000 ;
    END
  END PRDATA[1]
  PIN PRDATA[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 20.4375 47.8800 20.5125 48.3000 ;
    END
  END PRDATA[0]
  PIN PREADY
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.8625 0.0000 0.9375 0.5100 ;
    END
  END PREADY
  PIN PSLVERR
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 48.8400 47.3625 49.3500 47.4375 ;
    END
  END PSLVERR
  PIN pad_cfg_o[191]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 48.8400 22.7625 49.3500 22.8375 ;
    END
  END pad_cfg_o[191]
  PIN pad_cfg_o[190]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 18.5625 0.5100 18.6375 ;
    END
  END pad_cfg_o[190]
  PIN pad_cfg_o[189]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 48.8400 20.5125 49.3500 20.5875 ;
    END
  END pad_cfg_o[189]
  PIN pad_cfg_o[188]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 33.7125 0.5100 33.7875 ;
    END
  END pad_cfg_o[188]
  PIN pad_cfg_o[187]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 30.7125 47.7900 30.7875 48.3000 ;
    END
  END pad_cfg_o[187]
  PIN pad_cfg_o[186]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 48.8400 6.1125 49.3500 6.1875 ;
    END
  END pad_cfg_o[186]
  PIN pad_cfg_o[185]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 48.8400 28.7625 49.3500 28.8375 ;
    END
  END pad_cfg_o[185]
  PIN pad_cfg_o[184]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 48.8400 41.8125 49.3500 41.8875 ;
    END
  END pad_cfg_o[184]
  PIN pad_cfg_o[183]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 20.5125 0.5100 20.5875 ;
    END
  END pad_cfg_o[183]
  PIN pad_cfg_o[182]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9.0975 0.0000 9.1725 0.4200 ;
    END
  END pad_cfg_o[182]
  PIN pad_cfg_o[181]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 25.4625 0.0000 25.5375 0.5100 ;
    END
  END pad_cfg_o[181]
  PIN pad_cfg_o[180]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 38.4975 47.8800 38.5725 48.3000 ;
    END
  END pad_cfg_o[180]
  PIN pad_cfg_o[179]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 46.0575 0.0000 46.1325 0.4200 ;
    END
  END pad_cfg_o[179]
  PIN pad_cfg_o[178]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 25.4625 0.0000 25.5375 0.5100 ;
    END
  END pad_cfg_o[178]
  PIN pad_cfg_o[177]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 48.8400 12.8625 49.3500 12.9375 ;
    END
  END pad_cfg_o[177]
  PIN pad_cfg_o[176]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 48.8400 35.8125 49.3500 35.8875 ;
    END
  END pad_cfg_o[176]
  PIN pad_cfg_o[175]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18.7575 0.0000 18.8325 0.4200 ;
    END
  END pad_cfg_o[175]
  PIN pad_cfg_o[174]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 32.2125 47.7900 32.2875 48.3000 ;
    END
  END pad_cfg_o[174]
  PIN pad_cfg_o[173]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 25.2675 47.8800 25.3425 48.3000 ;
    END
  END pad_cfg_o[173]
  PIN pad_cfg_o[172]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10.7775 0.0000 10.8525 0.4200 ;
    END
  END pad_cfg_o[172]
  PIN pad_cfg_o[171]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 28.4625 0.0000 28.5375 0.5100 ;
    END
  END pad_cfg_o[171]
  PIN pad_cfg_o[170]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 19.1775 47.8800 19.2525 48.3000 ;
    END
  END pad_cfg_o[170]
  PIN pad_cfg_o[169]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 39.7125 0.5100 39.7875 ;
    END
  END pad_cfg_o[169]
  PIN pad_cfg_o[168]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 22.9125 47.7900 22.9875 48.3000 ;
    END
  END pad_cfg_o[168]
  PIN pad_cfg_o[167]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 48.8400 19.3125 49.3500 19.3875 ;
    END
  END pad_cfg_o[167]
  PIN pad_cfg_o[166]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 18.8625 0.5100 18.9375 ;
    END
  END pad_cfg_o[166]
  PIN pad_cfg_o[165]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 48.8400 20.3625 49.3500 20.4375 ;
    END
  END pad_cfg_o[165]
  PIN pad_cfg_o[164]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 31.0125 0.5100 31.0875 ;
    END
  END pad_cfg_o[164]
  PIN pad_cfg_o[163]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 48.8400 27.2625 49.3500 27.3375 ;
    END
  END pad_cfg_o[163]
  PIN pad_cfg_o[162]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 42.4875 0.0000 42.5625 0.4200 ;
    END
  END pad_cfg_o[162]
  PIN pad_cfg_o[161]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 48.8400 25.9125 49.3500 25.9875 ;
    END
  END pad_cfg_o[161]
  PIN pad_cfg_o[160]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 48.8400 39.4125 49.3500 39.4875 ;
    END
  END pad_cfg_o[160]
  PIN pad_cfg_o[159]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 21.2625 0.5100 21.3375 ;
    END
  END pad_cfg_o[159]
  PIN pad_cfg_o[158]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6.9975 0.0000 7.0725 0.4200 ;
    END
  END pad_cfg_o[158]
  PIN pad_cfg_o[157]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 22.3275 0.0000 22.4025 0.4200 ;
    END
  END pad_cfg_o[157]
  PIN pad_cfg_o[156]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 48.8400 38.5125 49.3500 38.5875 ;
    END
  END pad_cfg_o[156]
  PIN pad_cfg_o[155]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 42.4125 0.0000 42.4875 0.5100 ;
    END
  END pad_cfg_o[155]
  PIN pad_cfg_o[154]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 23.3625 0.0000 23.4375 0.5100 ;
    END
  END pad_cfg_o[154]
  PIN pad_cfg_o[153]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 48.8400 16.7625 49.3500 16.8375 ;
    END
  END pad_cfg_o[153]
  PIN pad_cfg_o[152]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 48.8400 32.8125 49.3500 32.8875 ;
    END
  END pad_cfg_o[152]
  PIN pad_cfg_o[151]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15.6075 0.0000 15.6825 0.4200 ;
    END
  END pad_cfg_o[151]
  PIN pad_cfg_o[150]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 31.9875 47.8800 32.0625 48.3000 ;
    END
  END pad_cfg_o[150]
  PIN pad_cfg_o[149]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 23.5875 47.8800 23.6625 48.3000 ;
    END
  END pad_cfg_o[149]
  PIN pad_cfg_o[148]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 7.6125 0.5100 7.6875 ;
    END
  END pad_cfg_o[148]
  PIN pad_cfg_o[147]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 31.3125 0.0000 31.3875 0.5100 ;
    END
  END pad_cfg_o[147]
  PIN pad_cfg_o[146]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 32.9625 0.5100 33.0375 ;
    END
  END pad_cfg_o[146]
  PIN pad_cfg_o[145]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 38.5125 0.5100 38.5875 ;
    END
  END pad_cfg_o[145]
  PIN pad_cfg_o[144]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 20.0175 47.8800 20.0925 48.3000 ;
    END
  END pad_cfg_o[144]
  PIN pad_cfg_o[143]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 48.8400 21.8625 49.3500 21.9375 ;
    END
  END pad_cfg_o[143]
  PIN pad_cfg_o[142]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 0.0000 16.5000 2.1225 17.1000 ;
    END
  END pad_cfg_o[142]
  PIN pad_cfg_o[141]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 29.8875 0.0000 29.9625 0.4200 ;
    END
  END pad_cfg_o[141]
  PIN pad_cfg_o[140]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 34.1625 0.5100 34.2375 ;
    END
  END pad_cfg_o[140]
  PIN pad_cfg_o[139]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 31.7625 47.7900 31.8375 48.3000 ;
    END
  END pad_cfg_o[139]
  PIN pad_cfg_o[138]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 48.8400 7.6125 49.3500 7.6875 ;
    END
  END pad_cfg_o[138]
  PIN pad_cfg_o[137]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 48.8400 27.8625 49.3500 27.9375 ;
    END
  END pad_cfg_o[137]
  PIN pad_cfg_o[136]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 48.8400 43.3125 49.3500 43.3875 ;
    END
  END pad_cfg_o[136]
  PIN pad_cfg_o[135]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 19.6125 0.5100 19.6875 ;
    END
  END pad_cfg_o[135]
  PIN pad_cfg_o[134]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9.7275 0.0000 9.8025 0.4200 ;
    END
  END pad_cfg_o[134]
  PIN pad_cfg_o[133]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 24.2175 0.0000 24.2925 0.4200 ;
    END
  END pad_cfg_o[133]
  PIN pad_cfg_o[132]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 37.3125 47.7900 37.3875 48.3000 ;
    END
  END pad_cfg_o[132]
  PIN pad_cfg_o[131]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 45.6375 0.0000 45.7125 0.4200 ;
    END
  END pad_cfg_o[131]
  PIN pad_cfg_o[130]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 24.2625 0.0000 24.3375 0.5100 ;
    END
  END pad_cfg_o[130]
  PIN pad_cfg_o[129]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 48.8400 13.6125 49.3500 13.6875 ;
    END
  END pad_cfg_o[129]
  PIN pad_cfg_o[128]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 48.8400 34.3125 49.3500 34.3875 ;
    END
  END pad_cfg_o[128]
  PIN pad_cfg_o[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17.8125 0.0000 17.8875 0.5100 ;
    END
  END pad_cfg_o[127]
  PIN pad_cfg_o[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 30.9375 47.8800 31.0125 48.3000 ;
    END
  END pad_cfg_o[126]
  PIN pad_cfg_o[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 24.2625 47.7900 24.3375 48.3000 ;
    END
  END pad_cfg_o[125]
  PIN pad_cfg_o[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11.1975 0.0000 11.2725 0.4200 ;
    END
  END pad_cfg_o[124]
  PIN pad_cfg_o[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 28.4625 0.0000 28.5375 0.5100 ;
    END
  END pad_cfg_o[123]
  PIN pad_cfg_o[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18.8625 47.7900 18.9375 48.3000 ;
    END
  END pad_cfg_o[122]
  PIN pad_cfg_o[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10.1475 47.8800 10.2225 48.3000 ;
    END
  END pad_cfg_o[121]
  PIN pad_cfg_o[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 22.5375 47.8800 22.6125 48.3000 ;
    END
  END pad_cfg_o[120]
  PIN pad_cfg_o[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 48.8400 22.1625 49.3500 22.2375 ;
    END
  END pad_cfg_o[119]
  PIN pad_cfg_o[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 14.8125 0.5100 14.8875 ;
    END
  END pad_cfg_o[118]
  PIN pad_cfg_o[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 27.5775 0.0000 27.6525 0.4200 ;
    END
  END pad_cfg_o[117]
  PIN pad_cfg_o[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 31.3125 0.5100 31.3875 ;
    END
  END pad_cfg_o[116]
  PIN pad_cfg_o[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 48.8400 27.5625 49.3500 27.6375 ;
    END
  END pad_cfg_o[115]
  PIN pad_cfg_o[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 41.2275 0.0000 41.3025 0.4200 ;
    END
  END pad_cfg_o[114]
  PIN pad_cfg_o[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 48.8400 25.6125 49.3500 25.6875 ;
    END
  END pad_cfg_o[113]
  PIN pad_cfg_o[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 43.5375 47.8800 43.6125 48.3000 ;
    END
  END pad_cfg_o[112]
  PIN pad_cfg_o[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18.8625 0.0000 18.9375 0.5100 ;
    END
  END pad_cfg_o[111]
  PIN pad_cfg_o[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10.7625 0.0000 10.8375 0.5100 ;
    END
  END pad_cfg_o[110]
  PIN pad_cfg_o[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 25.1625 0.0000 25.2375 0.5100 ;
    END
  END pad_cfg_o[109]
  PIN pad_cfg_o[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 40.5975 47.8800 40.6725 48.3000 ;
    END
  END pad_cfg_o[108]
  PIN pad_cfg_o[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 39.9675 0.0000 40.0425 0.4200 ;
    END
  END pad_cfg_o[107]
  PIN pad_cfg_o[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 25.1625 0.0000 25.2375 0.5100 ;
    END
  END pad_cfg_o[106]
  PIN pad_cfg_o[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 48.8400 13.0125 49.3500 13.0875 ;
    END
  END pad_cfg_o[105]
  PIN pad_cfg_o[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 48.8400 34.6125 49.3500 34.6875 ;
    END
  END pad_cfg_o[104]
  PIN pad_cfg_o[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 18.7125 0.0000 18.7875 0.5100 ;
    END
  END pad_cfg_o[103]
  PIN pad_cfg_o[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 28.3125 47.7900 28.3875 48.3000 ;
    END
  END pad_cfg_o[102]
  PIN pad_cfg_o[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 25.1625 47.7900 25.2375 48.3000 ;
    END
  END pad_cfg_o[101]
  PIN pad_cfg_o[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 11.2125 0.5100 11.2875 ;
    END
  END pad_cfg_o[100]
  PIN pad_cfg_o[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 32.0625 0.0000 32.1375 0.5100 ;
    END
  END pad_cfg_o[99]
  PIN pad_cfg_o[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18.5625 47.7900 18.6375 48.3000 ;
    END
  END pad_cfg_o[98]
  PIN pad_cfg_o[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 36.8625 0.5100 36.9375 ;
    END
  END pad_cfg_o[97]
  PIN pad_cfg_o[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17.9175 47.8800 17.9925 48.3000 ;
    END
  END pad_cfg_o[96]
  PIN pad_cfg_o[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 48.8400 18.8625 49.3500 18.9375 ;
    END
  END pad_cfg_o[95]
  PIN pad_cfg_o[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 22.9125 0.5100 22.9875 ;
    END
  END pad_cfg_o[94]
  PIN pad_cfg_o[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 48.8400 22.1625 49.3500 22.2375 ;
    END
  END pad_cfg_o[93]
  PIN pad_cfg_o[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 31.6125 0.5100 31.6875 ;
    END
  END pad_cfg_o[92]
  PIN pad_cfg_o[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 48.8400 31.0125 49.3500 31.0875 ;
    END
  END pad_cfg_o[91]
  PIN pad_cfg_o[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 48.8400 9.7125 49.3500 9.7875 ;
    END
  END pad_cfg_o[90]
  PIN pad_cfg_o[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 48.8400 26.0625 49.3500 26.1375 ;
    END
  END pad_cfg_o[89]
  PIN pad_cfg_o[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 48.8400 39.7125 49.3500 39.7875 ;
    END
  END pad_cfg_o[88]
  PIN pad_cfg_o[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 22.4625 0.5100 22.5375 ;
    END
  END pad_cfg_o[87]
  PIN pad_cfg_o[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5.9475 0.0000 6.0225 0.4200 ;
    END
  END pad_cfg_o[86]
  PIN pad_cfg_o[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 24.1125 0.0000 24.1875 0.5100 ;
    END
  END pad_cfg_o[85]
  PIN pad_cfg_o[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 37.4625 47.7900 37.5375 48.3000 ;
    END
  END pad_cfg_o[84]
  PIN pad_cfg_o[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 37.9125 0.0000 37.9875 0.5100 ;
    END
  END pad_cfg_o[83]
  PIN pad_cfg_o[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 21.8625 0.0000 21.9375 0.5100 ;
    END
  END pad_cfg_o[82]
  PIN pad_cfg_o[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 48.8400 15.5625 49.3500 15.6375 ;
    END
  END pad_cfg_o[81]
  PIN pad_cfg_o[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 48.8400 32.2125 49.3500 32.2875 ;
    END
  END pad_cfg_o[80]
  PIN pad_cfg_o[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16.6125 0.0000 16.6875 0.5100 ;
    END
  END pad_cfg_o[79]
  PIN pad_cfg_o[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 27.8625 47.7900 27.9375 48.3000 ;
    END
  END pad_cfg_o[78]
  PIN pad_cfg_o[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 25.3125 47.7900 25.3875 48.3000 ;
    END
  END pad_cfg_o[77]
  PIN pad_cfg_o[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 12.5625 0.5100 12.6375 ;
    END
  END pad_cfg_o[76]
  PIN pad_cfg_o[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 31.7625 0.0000 31.8375 0.5100 ;
    END
  END pad_cfg_o[75]
  PIN pad_cfg_o[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 31.1625 0.5100 31.2375 ;
    END
  END pad_cfg_o[74]
  PIN pad_cfg_o[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 37.1625 0.5100 37.2375 ;
    END
  END pad_cfg_o[73]
  PIN pad_cfg_o[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 22.1175 47.8800 22.1925 48.3000 ;
    END
  END pad_cfg_o[72]
  PIN pad_cfg_o[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 48.8400 20.0625 49.3500 20.1375 ;
    END
  END pad_cfg_o[71]
  PIN pad_cfg_o[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 20.2125 0.5100 20.2875 ;
    END
  END pad_cfg_o[70]
  PIN pad_cfg_o[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 48.8400 22.7625 49.3500 22.8375 ;
    END
  END pad_cfg_o[69]
  PIN pad_cfg_o[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 33.7125 0.5100 33.7875 ;
    END
  END pad_cfg_o[68]
  PIN pad_cfg_o[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 28.8375 47.8800 28.9125 48.3000 ;
    END
  END pad_cfg_o[67]
  PIN pad_cfg_o[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 48.8400 6.4125 49.3500 6.4875 ;
    END
  END pad_cfg_o[66]
  PIN pad_cfg_o[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 48.8400 28.9125 49.3500 28.9875 ;
    END
  END pad_cfg_o[65]
  PIN pad_cfg_o[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 48.8400 37.9125 49.3500 37.9875 ;
    END
  END pad_cfg_o[64]
  PIN pad_cfg_o[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 20.0625 0.5100 20.1375 ;
    END
  END pad_cfg_o[63]
  PIN pad_cfg_o[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5.6625 0.0000 5.7375 0.5100 ;
    END
  END pad_cfg_o[62]
  PIN pad_cfg_o[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 21.8625 0.5100 21.9375 ;
    END
  END pad_cfg_o[61]
  PIN pad_cfg_o[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 48.8400 37.3125 49.3500 37.3875 ;
    END
  END pad_cfg_o[60]
  PIN pad_cfg_o[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 41.2125 0.0000 41.2875 0.5100 ;
    END
  END pad_cfg_o[59]
  PIN pad_cfg_o[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 22.4625 0.0000 22.5375 0.5100 ;
    END
  END pad_cfg_o[58]
  PIN pad_cfg_o[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 48.8400 16.7625 49.3500 16.8375 ;
    END
  END pad_cfg_o[57]
  PIN pad_cfg_o[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 48.8400 31.9125 49.3500 31.9875 ;
    END
  END pad_cfg_o[56]
  PIN pad_cfg_o[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15.7125 0.0000 15.7875 0.5100 ;
    END
  END pad_cfg_o[55]
  PIN pad_cfg_o[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 31.5675 47.8800 31.6425 48.3000 ;
    END
  END pad_cfg_o[54]
  PIN pad_cfg_o[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 22.3125 47.7900 22.3875 48.3000 ;
    END
  END pad_cfg_o[53]
  PIN pad_cfg_o[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 8.9625 0.5100 9.0375 ;
    END
  END pad_cfg_o[52]
  PIN pad_cfg_o[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 32.5125 0.0000 32.5875 0.5100 ;
    END
  END pad_cfg_o[51]
  PIN pad_cfg_o[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 0.0000 33.3000 2.1225 33.9000 ;
    END
  END pad_cfg_o[50]
  PIN pad_cfg_o[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 36.8625 0.5100 36.9375 ;
    END
  END pad_cfg_o[49]
  PIN pad_cfg_o[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 19.4625 47.7900 19.5375 48.3000 ;
    END
  END pad_cfg_o[48]
  PIN pad_cfg_o[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 48.8400 23.0625 49.3500 23.1375 ;
    END
  END pad_cfg_o[47]
  PIN pad_cfg_o[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 14.2125 0.5100 14.2875 ;
    END
  END pad_cfg_o[46]
  PIN pad_cfg_o[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 28.2075 0.0000 28.2825 0.4200 ;
    END
  END pad_cfg_o[45]
  PIN pad_cfg_o[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 29.8125 0.5100 29.8875 ;
    END
  END pad_cfg_o[44]
  PIN pad_cfg_o[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 29.2575 47.8800 29.3325 48.3000 ;
    END
  END pad_cfg_o[43]
  PIN pad_cfg_o[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 48.8400 9.7125 49.3500 9.7875 ;
    END
  END pad_cfg_o[42]
  PIN pad_cfg_o[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 48.8400 27.2625 49.3500 27.3375 ;
    END
  END pad_cfg_o[41]
  PIN pad_cfg_o[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 42.4875 47.8800 42.5625 48.3000 ;
    END
  END pad_cfg_o[40]
  PIN pad_cfg_o[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 17.8125 0.0000 17.8875 0.5100 ;
    END
  END pad_cfg_o[39]
  PIN pad_cfg_o[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10.4625 0.0000 10.5375 0.5100 ;
    END
  END pad_cfg_o[38]
  PIN pad_cfg_o[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 25.8975 0.0000 25.9725 0.4200 ;
    END
  END pad_cfg_o[37]
  PIN pad_cfg_o[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 41.0625 47.7900 41.1375 48.3000 ;
    END
  END pad_cfg_o[36]
  PIN pad_cfg_o[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 38.7075 0.0000 38.7825 0.4200 ;
    END
  END pad_cfg_o[35]
  PIN pad_cfg_o[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 24.8625 0.0000 24.9375 0.5100 ;
    END
  END pad_cfg_o[34]
  PIN pad_cfg_o[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 48.8400 13.7625 49.3500 13.8375 ;
    END
  END pad_cfg_o[33]
  PIN pad_cfg_o[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 48.8400 33.8625 49.3500 33.9375 ;
    END
  END pad_cfg_o[32]
  PIN pad_cfg_o[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18.1125 0.0000 18.1875 0.5100 ;
    END
  END pad_cfg_o[31]
  PIN pad_cfg_o[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 27.1575 47.8800 27.2325 48.3000 ;
    END
  END pad_cfg_o[30]
  PIN pad_cfg_o[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 25.7625 47.7900 25.8375 48.3000 ;
    END
  END pad_cfg_o[29]
  PIN pad_cfg_o[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12.6675 0.0000 12.7425 0.4200 ;
    END
  END pad_cfg_o[28]
  PIN pad_cfg_o[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 29.6625 0.0000 29.7375 0.5100 ;
    END
  END pad_cfg_o[27]
  PIN pad_cfg_o[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 29.2125 0.5100 29.2875 ;
    END
  END pad_cfg_o[26]
  PIN pad_cfg_o[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10.9125 47.7900 10.9875 48.3000 ;
    END
  END pad_cfg_o[25]
  PIN pad_cfg_o[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15.8175 47.8800 15.8925 48.3000 ;
    END
  END pad_cfg_o[24]
  PIN pad_cfg_o[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 48.8400 19.6125 49.3500 19.6875 ;
    END
  END pad_cfg_o[23]
  PIN pad_cfg_o[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 23.2125 0.5100 23.2875 ;
    END
  END pad_cfg_o[22]
  PIN pad_cfg_o[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 48.8400 23.0625 49.3500 23.1375 ;
    END
  END pad_cfg_o[21]
  PIN pad_cfg_o[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 32.6625 0.5100 32.7375 ;
    END
  END pad_cfg_o[20]
  PIN pad_cfg_o[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 32.2125 47.7900 32.2875 48.3000 ;
    END
  END pad_cfg_o[19]
  PIN pad_cfg_o[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 48.8400 10.6125 49.3500 10.6875 ;
    END
  END pad_cfg_o[18]
  PIN pad_cfg_o[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 48.8400 24.5625 49.3500 24.6375 ;
    END
  END pad_cfg_o[17]
  PIN pad_cfg_o[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 48.8400 38.6625 49.3500 38.7375 ;
    END
  END pad_cfg_o[16]
  PIN pad_cfg_o[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 22.9125 0.5100 22.9875 ;
    END
  END pad_cfg_o[15]
  PIN pad_cfg_o[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7.4175 0.0000 7.4925 0.4200 ;
    END
  END pad_cfg_o[14]
  PIN pad_cfg_o[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 23.8125 0.0000 23.8875 0.5100 ;
    END
  END pad_cfg_o[13]
  PIN pad_cfg_o[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 48.8400 37.9125 49.3500 37.9875 ;
    END
  END pad_cfg_o[12]
  PIN pad_cfg_o[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 38.8125 0.0000 38.8875 0.5100 ;
    END
  END pad_cfg_o[11]
  PIN pad_cfg_o[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 21.2625 0.0000 21.3375 0.5100 ;
    END
  END pad_cfg_o[10]
  PIN pad_cfg_o[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 48.8400 16.3125 49.3500 16.3875 ;
    END
  END pad_cfg_o[9]
  PIN pad_cfg_o[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 48.8400 31.6125 49.3500 31.6875 ;
    END
  END pad_cfg_o[8]
  PIN pad_cfg_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16.0275 0.0000 16.1025 0.4200 ;
    END
  END pad_cfg_o[7]
  PIN pad_cfg_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 28.9125 47.7900 28.9875 48.3000 ;
    END
  END pad_cfg_o[6]
  PIN pad_cfg_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 23.9625 47.7900 24.0375 48.3000 ;
    END
  END pad_cfg_o[5]
  PIN pad_cfg_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 13.3125 0.5100 13.3875 ;
    END
  END pad_cfg_o[4]
  PIN pad_cfg_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 31.9125 0.0000 31.9875 0.5100 ;
    END
  END pad_cfg_o[3]
  PIN pad_cfg_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17.6625 47.7900 17.7375 48.3000 ;
    END
  END pad_cfg_o[2]
  PIN pad_cfg_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 36.4125 0.5100 36.4875 ;
    END
  END pad_cfg_o[1]
  PIN pad_cfg_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 21.6975 47.8800 21.7725 48.3000 ;
    END
  END pad_cfg_o[0]
  PIN clk_gate_o[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 23.9625 47.7900 24.0375 48.3000 ;
    END
  END clk_gate_o[31]
  PIN clk_gate_o[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 28.4625 0.5100 28.5375 ;
    END
  END clk_gate_o[30]
  PIN clk_gate_o[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 48.8400 19.4625 49.3500 19.5375 ;
    END
  END clk_gate_o[29]
  PIN clk_gate_o[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 19.4625 0.5100 19.5375 ;
    END
  END clk_gate_o[28]
  PIN clk_gate_o[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 31.9875 0.0000 32.0625 0.4200 ;
    END
  END clk_gate_o[27]
  PIN clk_gate_o[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 25.3125 0.5100 25.3875 ;
    END
  END clk_gate_o[26]
  PIN clk_gate_o[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 48.8400 24.8625 49.3500 24.9375 ;
    END
  END clk_gate_o[25]
  PIN clk_gate_o[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 36.8175 0.0000 36.8925 0.4200 ;
    END
  END clk_gate_o[24]
  PIN clk_gate_o[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 34.7625 0.5100 34.8375 ;
    END
  END clk_gate_o[23]
  PIN clk_gate_o[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 16.7625 0.5100 16.8375 ;
    END
  END clk_gate_o[22]
  PIN clk_gate_o[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 48.8400 25.1625 49.3500 25.2375 ;
    END
  END clk_gate_o[21]
  PIN clk_gate_o[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 33.6675 47.8800 33.7425 48.3000 ;
    END
  END clk_gate_o[20]
  PIN clk_gate_o[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15.1875 0.0000 15.2625 0.4200 ;
    END
  END clk_gate_o[19]
  PIN clk_gate_o[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 9.4125 0.5100 9.4875 ;
    END
  END clk_gate_o[18]
  PIN clk_gate_o[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 21.6975 0.0000 21.7725 0.4200 ;
    END
  END clk_gate_o[17]
  PIN clk_gate_o[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 37.7625 47.7900 37.8375 48.3000 ;
    END
  END clk_gate_o[16]
  PIN clk_gate_o[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3.6375 47.8800 3.7125 48.3000 ;
    END
  END clk_gate_o[15]
  PIN clk_gate_o[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 24.2625 0.5100 24.3375 ;
    END
  END clk_gate_o[14]
  PIN clk_gate_o[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 33.0375 0.0000 33.1125 0.4200 ;
    END
  END clk_gate_o[13]
  PIN clk_gate_o[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 22.7475 0.0000 22.8225 0.4200 ;
    END
  END clk_gate_o[12]
  PIN clk_gate_o[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 48.8400 16.1625 49.3500 16.2375 ;
    END
  END clk_gate_o[11]
  PIN clk_gate_o[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 48.8400 34.6125 49.3500 34.6875 ;
    END
  END clk_gate_o[10]
  PIN clk_gate_o[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18.1275 0.0000 18.2025 0.4200 ;
    END
  END clk_gate_o[9]
  PIN clk_gate_o[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 30.5175 47.8800 30.5925 48.3000 ;
    END
  END clk_gate_o[8]
  PIN clk_gate_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 46.0125 0.5100 46.0875 ;
    END
  END clk_gate_o[7]
  PIN clk_gate_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 22.4625 0.5100 22.5375 ;
    END
  END clk_gate_o[6]
  PIN clk_gate_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 25.4625 0.5100 25.5375 ;
    END
  END clk_gate_o[5]
  PIN clk_gate_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 11.9625 0.5100 12.0375 ;
    END
  END clk_gate_o[4]
  PIN clk_gate_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 29.0475 0.0000 29.1225 0.4200 ;
    END
  END clk_gate_o[3]
  PIN clk_gate_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 26.0625 0.5100 26.1375 ;
    END
  END clk_gate_o[2]
  PIN clk_gate_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9.5175 47.8800 9.5925 48.3000 ;
    END
  END clk_gate_o[1]
  PIN clk_gate_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 21.2775 47.8800 21.3525 48.3000 ;
    END
  END clk_gate_o[0]
  PIN pad_mux_o[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 25.4625 47.7900 25.5375 48.3000 ;
    END
  END pad_mux_o[31]
  PIN pad_mux_o[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 27.1125 0.5100 27.1875 ;
    END
  END pad_mux_o[30]
  PIN pad_mux_o[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 48.8400 21.4125 49.3500 21.4875 ;
    END
  END pad_mux_o[29]
  PIN pad_mux_o[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 15.2625 0.5100 15.3375 ;
    END
  END pad_mux_o[28]
  PIN pad_mux_o[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 31.6125 0.0000 31.6875 0.5100 ;
    END
  END pad_mux_o[27]
  PIN pad_mux_o[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 27.2625 0.5100 27.3375 ;
    END
  END pad_mux_o[26]
  PIN pad_mux_o[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 48.8400 26.5125 49.3500 26.5875 ;
    END
  END pad_mux_o[25]
  PIN pad_mux_o[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 37.4625 0.0000 37.5375 0.5100 ;
    END
  END pad_mux_o[24]
  PIN pad_mux_o[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 32.2125 0.5100 32.2875 ;
    END
  END pad_mux_o[23]
  PIN pad_mux_o[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 17.6625 0.5100 17.7375 ;
    END
  END pad_mux_o[22]
  PIN pad_mux_o[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 48.8400 26.5125 49.3500 26.5875 ;
    END
  END pad_mux_o[21]
  PIN pad_mux_o[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 35.5575 47.8800 35.6325 48.3000 ;
    END
  END pad_mux_o[20]
  PIN pad_mux_o[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16.1625 0.0000 16.2375 0.5100 ;
    END
  END pad_mux_o[19]
  PIN pad_mux_o[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 7.9125 0.5100 7.9875 ;
    END
  END pad_mux_o[18]
  PIN pad_mux_o[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 22.6125 0.0000 22.6875 0.5100 ;
    END
  END pad_mux_o[17]
  PIN pad_mux_o[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 36.1875 47.8800 36.2625 48.3000 ;
    END
  END pad_mux_o[16]
  PIN pad_mux_o[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 42.8625 0.5100 42.9375 ;
    END
  END pad_mux_o[15]
  PIN pad_mux_o[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 26.5125 0.5100 26.5875 ;
    END
  END pad_mux_o[14]
  PIN pad_mux_o[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 33.6675 0.0000 33.7425 0.4200 ;
    END
  END pad_mux_o[13]
  PIN pad_mux_o[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 23.9625 0.0000 24.0375 0.5100 ;
    END
  END pad_mux_o[12]
  PIN pad_mux_o[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 48.8400 15.1125 49.3500 15.1875 ;
    END
  END pad_mux_o[11]
  PIN pad_mux_o[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 48.8400 32.9625 49.3500 33.0375 ;
    END
  END pad_mux_o[10]
  PIN pad_mux_o[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 19.0125 0.0000 19.0875 0.5100 ;
    END
  END pad_mux_o[9]
  PIN pad_mux_o[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 31.0125 47.7900 31.0875 48.3000 ;
    END
  END pad_mux_o[8]
  PIN pad_mux_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 41.0625 0.5100 41.1375 ;
    END
  END pad_mux_o[7]
  PIN pad_mux_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 20.3625 0.5100 20.4375 ;
    END
  END pad_mux_o[6]
  PIN pad_mux_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 21.2625 47.7900 21.3375 48.3000 ;
    END
  END pad_mux_o[5]
  PIN pad_mux_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 13.3125 0.5100 13.3875 ;
    END
  END pad_mux_o[4]
  PIN pad_mux_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 29.0625 0.0000 29.1375 0.5100 ;
    END
  END pad_mux_o[3]
  PIN pad_mux_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 0.0000 26.1000 2.1225 26.7000 ;
    END
  END pad_mux_o[2]
  PIN pad_mux_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9.2625 47.7900 9.3375 48.3000 ;
    END
  END pad_mux_o[1]
  PIN pad_mux_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 19.9125 47.7900 19.9875 48.3000 ;
    END
  END pad_mux_o[0]
  PIN boot_addr_o[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 25.6875 47.8800 25.7625 48.3000 ;
    END
  END boot_addr_o[31]
  PIN boot_addr_o[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 26.3625 0.5100 26.4375 ;
    END
  END boot_addr_o[30]
  PIN boot_addr_o[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 48.8400 19.7625 49.3500 19.8375 ;
    END
  END boot_addr_o[29]
  PIN boot_addr_o[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 16.9125 0.5100 16.9875 ;
    END
  END boot_addr_o[28]
  PIN boot_addr_o[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 30.9375 0.0000 31.0125 0.4200 ;
    END
  END boot_addr_o[27]
  PIN boot_addr_o[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 26.8125 0.5100 26.8875 ;
    END
  END boot_addr_o[26]
  PIN boot_addr_o[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 48.8400 28.4625 49.3500 28.5375 ;
    END
  END boot_addr_o[25]
  PIN boot_addr_o[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 39.5475 0.0000 39.6225 0.4200 ;
    END
  END boot_addr_o[24]
  PIN boot_addr_o[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 33.2625 0.5100 33.3375 ;
    END
  END boot_addr_o[23]
  PIN boot_addr_o[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 17.9625 0.5100 18.0375 ;
    END
  END boot_addr_o[22]
  PIN boot_addr_o[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 48.8400 28.6125 49.3500 28.6875 ;
    END
  END boot_addr_o[21]
  PIN boot_addr_o[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 37.1625 47.7900 37.2375 48.3000 ;
    END
  END boot_addr_o[20]
  PIN boot_addr_o[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17.0625 0.0000 17.1375 0.5100 ;
    END
  END boot_addr_o[19]
  PIN boot_addr_o[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 7.1625 0.5100 7.2375 ;
    END
  END boot_addr_o[18]
  PIN boot_addr_o[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 23.6625 0.0000 23.7375 0.5100 ;
    END
  END boot_addr_o[17]
  PIN boot_addr_o[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 39.5475 47.8800 39.6225 48.3000 ;
    END
  END boot_addr_o[16]
  PIN boot_addr_o[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 43.6125 0.5100 43.6875 ;
    END
  END boot_addr_o[15]
  PIN boot_addr_o[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 26.6625 0.5100 26.7375 ;
    END
  END boot_addr_o[14]
  PIN boot_addr_o[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 37.7625 0.0000 37.8375 0.5100 ;
    END
  END boot_addr_o[13]
  PIN boot_addr_o[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 25.0575 0.0000 25.1325 0.4200 ;
    END
  END boot_addr_o[12]
  PIN boot_addr_o[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 48.8400 15.5625 49.3500 15.6375 ;
    END
  END boot_addr_o[11]
  PIN boot_addr_o[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 48.8400 31.9125 49.3500 31.9875 ;
    END
  END boot_addr_o[10]
  PIN boot_addr_o[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 17.2125 0.0000 17.2875 0.5100 ;
    END
  END boot_addr_o[9]
  PIN boot_addr_o[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 28.4175 47.8800 28.4925 48.3000 ;
    END
  END boot_addr_o[8]
  PIN boot_addr_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 40.4625 0.5100 40.5375 ;
    END
  END boot_addr_o[7]
  PIN boot_addr_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 22.0125 0.5100 22.0875 ;
    END
  END boot_addr_o[6]
  PIN boot_addr_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 24.2625 47.7900 24.3375 48.3000 ;
    END
  END boot_addr_o[5]
  PIN boot_addr_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 11.3625 0.5100 11.4375 ;
    END
  END boot_addr_o[4]
  PIN boot_addr_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 30.3075 0.0000 30.3825 0.4200 ;
    END
  END boot_addr_o[3]
  PIN boot_addr_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 29.6625 0.5100 29.7375 ;
    END
  END boot_addr_o[2]
  PIN boot_addr_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9.0975 47.8800 9.1725 48.3000 ;
    END
  END boot_addr_o[1]
  PIN boot_addr_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 23.1675 47.8800 23.2425 48.3000 ;
    END
  END boot_addr_o[0]
  OBS
    LAYER M1 ;
        RECT 0.0000 0.0000 49.3500 48.3000 ;
    LAYER M2 ;
        RECT 0.0000 0.0000 49.3500 48.3000 ;
    LAYER M3 ;
        RECT 0.0000 0.0000 49.3500 48.3000 ;
    LAYER M4 ;
        RECT 0.0000 0.0000 49.3500 48.3000 ;
    LAYER M5 ;
        RECT 0.0000 0.0000 49.3500 48.3000 ;
    LAYER M6 ;
        RECT 0.0000 0.0000 49.3500 48.3000 ;
    LAYER M7 ;
        RECT 0.0000 0.0000 49.3500 48.3000 ;
    LAYER M8 ;
        RECT 0.0000 0.0000 49.3500 48.3000 ;
  END
END apb_pulpino


VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO apb_spi_master
  CLASS BLOCK ;
    SIZE 88.4100 BY 88.2000 ;
  FOREIGN apb_spi_master 0.000000 0.000000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN HCLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 41.9625 0.5100 42.0375 ;
    END
  END HCLK
  PIN HRESETn
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 42.0675 0.0000 42.1425 0.4200 ;
    END
  END HRESETn
  PIN PADDR[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 44.1675 87.7800 44.2425 88.2000 ;
    END
  END PADDR[11]
  PIN PADDR[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 44.1675 0.0000 44.2425 0.4200 ;
    END
  END PADDR[10]
  PIN PADDR[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 44.2125 87.6900 44.2875 88.2000 ;
    END
  END PADDR[9]
  PIN PADDR[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 44.2125 87.6900 44.2875 88.2000 ;
    END
  END PADDR[8]
  PIN PADDR[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 44.2125 0.0000 44.2875 0.5100 ;
    END
  END PADDR[7]
  PIN PADDR[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 44.2125 0.0000 44.2875 0.5100 ;
    END
  END PADDR[6]
  PIN PADDR[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 87.9000 47.3625 88.4100 47.4375 ;
    END
  END PADDR[5]
  PIN PADDR[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 87.9000 46.1625 88.4100 46.2375 ;
    END
  END PADDR[4]
  PIN PADDR[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 87.9000 46.6125 88.4100 46.6875 ;
    END
  END PADDR[3]
  PIN PADDR[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 87.9000 45.4125 88.4100 45.4875 ;
    END
  END PADDR[2]
  PIN PADDR[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 44.0625 0.5100 44.1375 ;
    END
  END PADDR[1]
  PIN PADDR[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 44.0625 0.5100 44.1375 ;
    END
  END PADDR[0]
  PIN PWDATA[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 87.9000 33.1125 88.4100 33.1875 ;
    END
  END PWDATA[31]
  PIN PWDATA[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 55.7175 0.0000 55.7925 0.4200 ;
    END
  END PWDATA[30]
  PIN PWDATA[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 59.7075 0.0000 59.7825 0.4200 ;
    END
  END PWDATA[29]
  PIN PWDATA[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 46.8975 0.0000 46.9725 0.4200 ;
    END
  END PWDATA[28]
  PIN PWDATA[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 43.9125 0.0000 43.9875 0.5100 ;
    END
  END PWDATA[27]
  PIN PWDATA[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 51.3075 0.0000 51.3825 0.4200 ;
    END
  END PWDATA[26]
  PIN PWDATA[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 47.7375 0.0000 47.8125 0.4200 ;
    END
  END PWDATA[25]
  PIN PWDATA[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 50.4675 0.0000 50.5425 0.4200 ;
    END
  END PWDATA[24]
  PIN PWDATA[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 62.2275 0.0000 62.3025 0.4200 ;
    END
  END PWDATA[23]
  PIN PWDATA[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 61.1775 0.0000 61.2525 0.4200 ;
    END
  END PWDATA[22]
  PIN PWDATA[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 87.9000 26.2125 88.4100 26.2875 ;
    END
  END PWDATA[21]
  PIN PWDATA[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 20.4375 0.0000 20.5125 0.4200 ;
    END
  END PWDATA[20]
  PIN PWDATA[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 34.9125 0.0000 34.9875 0.5100 ;
    END
  END PWDATA[19]
  PIN PWDATA[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 22.6125 0.5100 22.6875 ;
    END
  END PWDATA[18]
  PIN PWDATA[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 38.2875 0.0000 38.3625 0.4200 ;
    END
  END PWDATA[17]
  PIN PWDATA[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 26.6625 0.5100 26.7375 ;
    END
  END PWDATA[16]
  PIN PWDATA[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 23.1675 0.0000 23.2425 0.4200 ;
    END
  END PWDATA[15]
  PIN PWDATA[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17.2875 0.0000 17.3625 0.4200 ;
    END
  END PWDATA[14]
  PIN PWDATA[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 67.2675 0.0000 67.3425 0.4200 ;
    END
  END PWDATA[13]
  PIN PWDATA[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 29.2575 0.0000 29.3325 0.4200 ;
    END
  END PWDATA[12]
  PIN PWDATA[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 31.1475 0.0000 31.2225 0.4200 ;
    END
  END PWDATA[11]
  PIN PWDATA[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 31.3125 0.0000 31.3875 0.5100 ;
    END
  END PWDATA[10]
  PIN PWDATA[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 34.3125 0.0000 34.3875 0.5100 ;
    END
  END PWDATA[9]
  PIN PWDATA[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 31.5675 0.0000 31.6425 0.4200 ;
    END
  END PWDATA[8]
  PIN PWDATA[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 87.9000 30.8625 88.4100 30.9375 ;
    END
  END PWDATA[7]
  PIN PWDATA[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 87.9000 27.2625 88.4100 27.3375 ;
    END
  END PWDATA[6]
  PIN PWDATA[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 87.9000 18.4125 88.4100 18.4875 ;
    END
  END PWDATA[5]
  PIN PWDATA[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 87.9000 23.6625 88.4100 23.7375 ;
    END
  END PWDATA[4]
  PIN PWDATA[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 87.9000 20.3625 88.4100 20.4375 ;
    END
  END PWDATA[3]
  PIN PWDATA[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 87.9000 32.5125 88.4100 32.5875 ;
    END
  END PWDATA[2]
  PIN PWDATA[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 87.9000 31.4625 88.4100 31.5375 ;
    END
  END PWDATA[1]
  PIN PWDATA[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 87.9000 33.4125 88.4100 33.4875 ;
    END
  END PWDATA[0]
  PIN PWRITE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 87.9000 49.0125 88.4100 49.0875 ;
    END
  END PWRITE
  PIN PSEL
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 87.9000 48.2625 88.4100 48.3375 ;
    END
  END PSEL
  PIN PENABLE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 87.9000 48.2625 88.4100 48.3375 ;
    END
  END PENABLE
  PIN PRDATA[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 87.9000 45.4125 88.4100 45.4875 ;
    END
  END PRDATA[31]
  PIN PRDATA[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 86.2875 45.3000 88.4100 45.9000 ;
    END
  END PRDATA[30]
  PIN PRDATA[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 87.9000 32.2125 88.4100 32.2875 ;
    END
  END PRDATA[29]
  PIN PRDATA[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 49.8375 87.7800 49.9125 88.2000 ;
    END
  END PRDATA[28]
  PIN PRDATA[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 46.8975 87.7800 46.9725 88.2000 ;
    END
  END PRDATA[27]
  PIN PRDATA[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 51.5175 87.7800 51.5925 88.2000 ;
    END
  END PRDATA[26]
  PIN PRDATA[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 48.3675 87.7800 48.4425 88.2000 ;
    END
  END PRDATA[25]
  PIN PRDATA[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 49.7625 87.6900 49.8375 88.2000 ;
    END
  END PRDATA[24]
  PIN PRDATA[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 87.9000 32.8125 88.4100 32.8875 ;
    END
  END PRDATA[23]
  PIN PRDATA[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 87.9000 34.3125 88.4100 34.3875 ;
    END
  END PRDATA[22]
  PIN PRDATA[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 87.9000 32.5125 88.4100 32.5875 ;
    END
  END PRDATA[21]
  PIN PRDATA[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 39.5475 87.7800 39.6225 88.2000 ;
    END
  END PRDATA[20]
  PIN PRDATA[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 38.4975 87.7800 38.5725 88.2000 ;
    END
  END PRDATA[19]
  PIN PRDATA[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 37.6575 87.7800 37.7325 88.2000 ;
    END
  END PRDATA[18]
  PIN PRDATA[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 39.9675 87.7800 40.0425 88.2000 ;
    END
  END PRDATA[17]
  PIN PRDATA[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 38.0775 87.7800 38.1525 88.2000 ;
    END
  END PRDATA[16]
  PIN PRDATA[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 34.2975 0.0000 34.3725 0.4200 ;
    END
  END PRDATA[15]
  PIN PRDATA[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 35.1375 0.0000 35.2125 0.4200 ;
    END
  END PRDATA[14]
  PIN PRDATA[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 87.9000 33.1125 88.4100 33.1875 ;
    END
  END PRDATA[13]
  PIN PRDATA[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 38.5125 0.5100 38.5875 ;
    END
  END PRDATA[12]
  PIN PRDATA[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 45.4125 0.5100 45.4875 ;
    END
  END PRDATA[11]
  PIN PRDATA[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 45.4125 0.5100 45.4875 ;
    END
  END PRDATA[10]
  PIN PRDATA[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 43.3125 0.5100 43.3875 ;
    END
  END PRDATA[9]
  PIN PRDATA[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 44.8125 0.5100 44.8875 ;
    END
  END PRDATA[8]
  PIN PRDATA[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 87.9000 37.0125 88.4100 37.0875 ;
    END
  END PRDATA[7]
  PIN PRDATA[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 87.9000 40.6125 88.4100 40.6875 ;
    END
  END PRDATA[6]
  PIN PRDATA[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 87.9000 45.8625 88.4100 45.9375 ;
    END
  END PRDATA[5]
  PIN PRDATA[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 87.9000 48.5625 88.4100 48.6375 ;
    END
  END PRDATA[4]
  PIN PRDATA[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 87.9000 47.9625 88.4100 48.0375 ;
    END
  END PRDATA[3]
  PIN PRDATA[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 87.9000 48.5625 88.4100 48.6375 ;
    END
  END PRDATA[2]
  PIN PRDATA[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 87.9000 46.4625 88.4100 46.5375 ;
    END
  END PRDATA[1]
  PIN PRDATA[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 87.9000 45.8625 88.4100 45.9375 ;
    END
  END PRDATA[0]
  PIN PREADY
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 87.5625 87.6900 87.6375 88.2000 ;
    END
  END PREADY
  PIN PSLVERR
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 87.5625 87.6900 87.6375 88.2000 ;
    END
  END PSLVERR
  PIN events_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 87.9000 63.7125 88.4100 63.7875 ;
    END
  END events_o[1]
  PIN events_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 46.6125 87.6900 46.6875 88.2000 ;
    END
  END events_o[0]
  PIN spi_clk
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 87.9000 66.8625 88.4100 66.9375 ;
    END
  END spi_clk
  PIN spi_csn0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 42.6975 87.7800 42.7725 88.2000 ;
    END
  END spi_csn0
  PIN spi_csn1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 43.7475 87.7800 43.8225 88.2000 ;
    END
  END spi_csn1
  PIN spi_csn2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 42.2775 87.7800 42.3525 88.2000 ;
    END
  END spi_csn2
  PIN spi_csn3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 41.6475 87.7800 41.7225 88.2000 ;
    END
  END spi_csn3
  PIN spi_mode[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 87.9000 68.9625 88.4100 69.0375 ;
    END
  END spi_mode[1]
  PIN spi_mode[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 87.9000 55.9125 88.4100 55.9875 ;
    END
  END spi_mode[0]
  PIN spi_sdo0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 87.9000 40.7625 88.4100 40.8375 ;
    END
  END spi_sdo0
  PIN spi_sdo1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 55.7625 0.0000 55.8375 0.5100 ;
    END
  END spi_sdo1
  PIN spi_sdo2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 87.9000 36.5625 88.4100 36.6375 ;
    END
  END spi_sdo2
  PIN spi_sdo3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 87.9000 38.8125 88.4100 38.8875 ;
    END
  END spi_sdo3
  PIN spi_sdi0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 22.3275 87.7800 22.4025 88.2000 ;
    END
  END spi_sdi0
  PIN spi_sdi1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 63.4125 0.5100 63.4875 ;
    END
  END spi_sdi1
  PIN spi_sdi2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 61.3125 0.5100 61.3875 ;
    END
  END spi_sdi2
  PIN spi_sdi3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 61.0125 0.5100 61.0875 ;
    END
  END spi_sdi3
  OBS
    LAYER M1 ;
        RECT 0.0000 0.0000 88.4100 88.2000 ;
    LAYER M2 ;
        RECT 0.0000 0.0000 88.4100 88.2000 ;
    LAYER M3 ;
        RECT 0.0000 0.0000 88.4100 88.2000 ;
    LAYER M4 ;
        RECT 0.0000 0.0000 88.4100 88.2000 ;
    LAYER M5 ;
        RECT 0.0000 0.0000 88.4100 88.2000 ;
    LAYER M6 ;
        RECT 0.0000 0.0000 88.4100 88.2000 ;
    LAYER M7 ;
        RECT 0.0000 0.0000 88.4100 88.2000 ;
    LAYER M8 ;
        RECT 0.0000 0.0000 88.4100 88.2000 ;
  END
END apb_spi_master


VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO apb_timer
  CLASS BLOCK ;
    SIZE 52.9200 BY 52.5000 ;
  FOREIGN apb_timer 0.000000 0.000000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN HCLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 25.8975 0.0000 25.9725 0.4200 ;
    END
  END HCLK
  PIN HRESETn
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 26.6625 0.0000 26.7375 0.5100 ;
    END
  END HRESETn
  PIN PADDR[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 26.3175 52.0800 26.3925 52.5000 ;
    END
  END PADDR[11]
  PIN PADDR[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 26.3625 51.9900 26.4375 52.5000 ;
    END
  END PADDR[10]
  PIN PADDR[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 26.3625 51.9900 26.4375 52.5000 ;
    END
  END PADDR[9]
  PIN PADDR[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 26.3175 0.0000 26.3925 0.4200 ;
    END
  END PADDR[8]
  PIN PADDR[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 26.3625 0.0000 26.4375 0.5100 ;
    END
  END PADDR[7]
  PIN PADDR[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 26.3625 0.0000 26.4375 0.5100 ;
    END
  END PADDR[6]
  PIN PADDR[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 26.2125 0.5100 26.2875 ;
    END
  END PADDR[5]
  PIN PADDR[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 52.4100 25.4625 52.9200 25.5375 ;
    END
  END PADDR[4]
  PIN PADDR[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 52.4100 26.0625 52.9200 26.1375 ;
    END
  END PADDR[3]
  PIN PADDR[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 52.4100 26.2125 52.9200 26.2875 ;
    END
  END PADDR[2]
  PIN PADDR[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 26.2125 0.5100 26.2875 ;
    END
  END PADDR[1]
  PIN PADDR[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 26.7375 52.0800 26.8125 52.5000 ;
    END
  END PADDR[0]
  PIN PWDATA[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 27.1125 0.5100 27.1875 ;
    END
  END PWDATA[31]
  PIN PWDATA[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 27.4125 0.5100 27.4875 ;
    END
  END PWDATA[30]
  PIN PWDATA[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 24.7125 0.5100 24.7875 ;
    END
  END PWDATA[29]
  PIN PWDATA[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 28.7625 0.5100 28.8375 ;
    END
  END PWDATA[28]
  PIN PWDATA[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 24.7125 0.5100 24.7875 ;
    END
  END PWDATA[27]
  PIN PWDATA[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 23.9625 0.5100 24.0375 ;
    END
  END PWDATA[26]
  PIN PWDATA[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 23.9625 0.5100 24.0375 ;
    END
  END PWDATA[25]
  PIN PWDATA[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 27.4125 0.5100 27.4875 ;
    END
  END PWDATA[24]
  PIN PWDATA[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 0.0000 23.7000 2.1225 24.3000 ;
    END
  END PWDATA[23]
  PIN PWDATA[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 23.6625 0.5100 23.7375 ;
    END
  END PWDATA[22]
  PIN PWDATA[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 27.7125 0.5100 27.7875 ;
    END
  END PWDATA[21]
  PIN PWDATA[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 27.7125 0.5100 27.7875 ;
    END
  END PWDATA[20]
  PIN PWDATA[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 28.0125 0.5100 28.0875 ;
    END
  END PWDATA[19]
  PIN PWDATA[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 23.6625 0.5100 23.7375 ;
    END
  END PWDATA[18]
  PIN PWDATA[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 24.6375 0.0000 24.7125 0.4200 ;
    END
  END PWDATA[17]
  PIN PWDATA[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 23.3625 0.5100 23.4375 ;
    END
  END PWDATA[16]
  PIN PWDATA[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 52.4100 27.2625 52.9200 27.3375 ;
    END
  END PWDATA[15]
  PIN PWDATA[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 52.4100 24.7125 52.9200 24.7875 ;
    END
  END PWDATA[14]
  PIN PWDATA[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 52.4100 27.4125 52.9200 27.4875 ;
    END
  END PWDATA[13]
  PIN PWDATA[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 52.4100 24.5625 52.9200 24.6375 ;
    END
  END PWDATA[12]
  PIN PWDATA[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 52.4100 23.9625 52.9200 24.0375 ;
    END
  END PWDATA[11]
  PIN PWDATA[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 52.4100 27.5625 52.9200 27.6375 ;
    END
  END PWDATA[10]
  PIN PWDATA[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 52.4100 23.9625 52.9200 24.0375 ;
    END
  END PWDATA[9]
  PIN PWDATA[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 52.4100 27.7125 52.9200 27.7875 ;
    END
  END PWDATA[8]
  PIN PWDATA[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 50.7975 23.7000 52.9200 24.3000 ;
    END
  END PWDATA[7]
  PIN PWDATA[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 52.4100 23.6625 52.9200 23.7375 ;
    END
  END PWDATA[6]
  PIN PWDATA[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 52.4100 27.8625 52.9200 27.9375 ;
    END
  END PWDATA[5]
  PIN PWDATA[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 52.4100 28.0125 52.9200 28.0875 ;
    END
  END PWDATA[4]
  PIN PWDATA[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 52.4100 28.1625 52.9200 28.2375 ;
    END
  END PWDATA[3]
  PIN PWDATA[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 52.4100 23.6625 52.9200 23.7375 ;
    END
  END PWDATA[2]
  PIN PWDATA[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 52.4100 28.3125 52.9200 28.3875 ;
    END
  END PWDATA[1]
  PIN PWDATA[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 27.7875 0.0000 27.8625 0.4200 ;
    END
  END PWDATA[0]
  PIN PWRITE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 52.4100 28.4625 52.9200 28.5375 ;
    END
  END PWRITE
  PIN PSEL
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 52.4100 23.3625 52.9200 23.4375 ;
    END
  END PSEL
  PIN PENABLE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 52.4100 28.6125 52.9200 28.6875 ;
    END
  END PENABLE
  PIN PRDATA[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 25.9125 0.5100 25.9875 ;
    END
  END PRDATA[31]
  PIN PRDATA[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 25.9125 0.5100 25.9875 ;
    END
  END PRDATA[30]
  PIN PRDATA[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 0.0000 26.1000 2.1225 26.7000 ;
    END
  END PRDATA[29]
  PIN PRDATA[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 25.6125 0.5100 25.6875 ;
    END
  END PRDATA[28]
  PIN PRDATA[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 26.5125 0.5100 26.5875 ;
    END
  END PRDATA[27]
  PIN PRDATA[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 25.6125 0.5100 25.6875 ;
    END
  END PRDATA[26]
  PIN PRDATA[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 26.5125 0.5100 26.5875 ;
    END
  END PRDATA[25]
  PIN PRDATA[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 26.8125 0.5100 26.8875 ;
    END
  END PRDATA[24]
  PIN PRDATA[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 25.3125 0.5100 25.3875 ;
    END
  END PRDATA[23]
  PIN PRDATA[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 25.3125 0.5100 25.3875 ;
    END
  END PRDATA[22]
  PIN PRDATA[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 24.2625 0.5100 24.3375 ;
    END
  END PRDATA[21]
  PIN PRDATA[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 26.8125 0.5100 26.8875 ;
    END
  END PRDATA[20]
  PIN PRDATA[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 25.0125 0.5100 25.0875 ;
    END
  END PRDATA[19]
  PIN PRDATA[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 24.2625 0.5100 24.3375 ;
    END
  END PRDATA[18]
  PIN PRDATA[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 27.1125 0.5100 27.1875 ;
    END
  END PRDATA[17]
  PIN PRDATA[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 25.0125 0.5100 25.0875 ;
    END
  END PRDATA[16]
  PIN PRDATA[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 52.4100 25.9125 52.9200 25.9875 ;
    END
  END PRDATA[15]
  PIN PRDATA[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 52.4100 25.7625 52.9200 25.8375 ;
    END
  END PRDATA[14]
  PIN PRDATA[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 52.4100 26.3625 52.9200 26.4375 ;
    END
  END PRDATA[13]
  PIN PRDATA[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 50.7975 26.1000 52.9200 26.7000 ;
    END
  END PRDATA[12]
  PIN PRDATA[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 52.4100 26.5125 52.9200 26.5875 ;
    END
  END PRDATA[11]
  PIN PRDATA[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 52.4100 26.6625 52.9200 26.7375 ;
    END
  END PRDATA[10]
  PIN PRDATA[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 52.4100 25.6125 52.9200 25.6875 ;
    END
  END PRDATA[9]
  PIN PRDATA[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 52.4100 25.3125 52.9200 25.3875 ;
    END
  END PRDATA[8]
  PIN PRDATA[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 52.4100 24.2625 52.9200 24.3375 ;
    END
  END PRDATA[7]
  PIN PRDATA[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 52.4100 26.8125 52.9200 26.8875 ;
    END
  END PRDATA[6]
  PIN PRDATA[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 52.4100 24.2625 52.9200 24.3375 ;
    END
  END PRDATA[5]
  PIN PRDATA[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 52.4100 25.1625 52.9200 25.2375 ;
    END
  END PRDATA[4]
  PIN PRDATA[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 52.4100 26.9625 52.9200 27.0375 ;
    END
  END PRDATA[3]
  PIN PRDATA[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 52.4100 25.0125 52.9200 25.0875 ;
    END
  END PRDATA[2]
  PIN PRDATA[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 52.4100 27.1125 52.9200 27.1875 ;
    END
  END PRDATA[1]
  PIN PRDATA[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 52.4100 24.8625 52.9200 24.9375 ;
    END
  END PRDATA[0]
  PIN PREADY
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 52.0125 0.0000 52.0875 0.5100 ;
    END
  END PREADY
  PIN PSLVERR
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 0.8625 0.5100 0.9375 ;
    END
  END PSLVERR
  PIN irq_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 26.7375 0.0000 26.8125 0.4200 ;
    END
  END irq_o[3]
  PIN irq_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 25.2675 0.0000 25.3425 0.4200 ;
    END
  END irq_o[2]
  PIN irq_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 26.8125 51.9900 26.8875 52.5000 ;
    END
  END irq_o[1]
  PIN irq_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 25.2675 52.0800 25.3425 52.5000 ;
    END
  END irq_o[0]
  OBS
    LAYER M1 ;
        RECT 0.0000 0.0000 52.9200 52.5000 ;
    LAYER M2 ;
        RECT 0.0000 0.0000 52.9200 52.5000 ;
    LAYER M3 ;
        RECT 0.0000 0.0000 52.9200 52.5000 ;
    LAYER M4 ;
        RECT 0.0000 0.0000 52.9200 52.5000 ;
    LAYER M5 ;
        RECT 0.0000 0.0000 52.9200 52.5000 ;
    LAYER M6 ;
        RECT 0.0000 0.0000 52.9200 52.5000 ;
    LAYER M7 ;
        RECT 0.0000 0.0000 52.9200 52.5000 ;
    LAYER M8 ;
        RECT 0.0000 0.0000 52.9200 52.5000 ;
  END
END apb_timer


VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO apb_uart
  CLASS BLOCK ;
    SIZE 110.4600 BY 110.2500 ;
  FOREIGN apb_uart 0.000000 0.000000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 54.6675 0.0000 54.7425 0.4200 ;
    END
  END CLK
  PIN RSTN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 109.9500 54.7125 110.4600 54.7875 ;
    END
  END RSTN
  PIN PSEL
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 63.4875 0.0000 63.5625 0.4200 ;
    END
  END PSEL
  PIN PENABLE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 63.5625 0.0000 63.6375 0.5100 ;
    END
  END PENABLE
  PIN PWRITE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 62.8575 0.0000 62.9325 0.4200 ;
    END
  END PWRITE
  PIN PADDR[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 73.9875 0.0000 74.0625 0.4200 ;
    END
  END PADDR[2]
  PIN PADDR[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 75.0375 0.0000 75.1125 0.4200 ;
    END
  END PADDR[1]
  PIN PADDR[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 74.6175 0.0000 74.6925 0.4200 ;
    END
  END PADDR[0]
  PIN PWDATA[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 55.0875 109.8300 55.1625 110.2500 ;
    END
  END PWDATA[31]
  PIN PWDATA[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 55.1625 109.7400 55.2375 110.2500 ;
    END
  END PWDATA[30]
  PIN PWDATA[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 55.1625 109.7400 55.2375 110.2500 ;
    END
  END PWDATA[29]
  PIN PWDATA[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 55.0875 0.0000 55.1625 0.4200 ;
    END
  END PWDATA[28]
  PIN PWDATA[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 55.1625 0.0000 55.2375 0.5100 ;
    END
  END PWDATA[27]
  PIN PWDATA[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 55.1625 0.0000 55.2375 0.5100 ;
    END
  END PWDATA[26]
  PIN PWDATA[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 55.0125 0.5100 55.0875 ;
    END
  END PWDATA[25]
  PIN PWDATA[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 55.0125 0.5100 55.0875 ;
    END
  END PWDATA[24]
  PIN PWDATA[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 0.0000 54.9000 2.1225 55.5000 ;
    END
  END PWDATA[23]
  PIN PWDATA[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 109.9500 55.0125 110.4600 55.0875 ;
    END
  END PWDATA[22]
  PIN PWDATA[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 109.9500 55.0125 110.4600 55.0875 ;
    END
  END PWDATA[21]
  PIN PWDATA[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 108.3375 54.9000 110.4600 55.5000 ;
    END
  END PWDATA[20]
  PIN PWDATA[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 55.5075 109.8300 55.5825 110.2500 ;
    END
  END PWDATA[19]
  PIN PWDATA[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 55.4625 109.7400 55.5375 110.2500 ;
    END
  END PWDATA[18]
  PIN PWDATA[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 55.4625 109.7400 55.5375 110.2500 ;
    END
  END PWDATA[17]
  PIN PWDATA[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 55.5075 0.0000 55.5825 0.4200 ;
    END
  END PWDATA[16]
  PIN PWDATA[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 55.4625 0.0000 55.5375 0.5100 ;
    END
  END PWDATA[15]
  PIN PWDATA[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 55.4625 0.0000 55.5375 0.5100 ;
    END
  END PWDATA[14]
  PIN PWDATA[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 55.3125 0.5100 55.3875 ;
    END
  END PWDATA[13]
  PIN PWDATA[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 55.3125 0.5100 55.3875 ;
    END
  END PWDATA[12]
  PIN PWDATA[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 54.8625 109.7400 54.9375 110.2500 ;
    END
  END PWDATA[11]
  PIN PWDATA[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 54.8625 109.7400 54.9375 110.2500 ;
    END
  END PWDATA[10]
  PIN PWDATA[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 109.9500 55.3125 110.4600 55.3875 ;
    END
  END PWDATA[9]
  PIN PWDATA[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 109.9500 55.3125 110.4600 55.3875 ;
    END
  END PWDATA[8]
  PIN PWDATA[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 109.9500 32.9625 110.4600 33.0375 ;
    END
  END PWDATA[7]
  PIN PWDATA[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 109.9500 25.7625 110.4600 25.8375 ;
    END
  END PWDATA[6]
  PIN PWDATA[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 109.9500 24.5625 110.4600 24.6375 ;
    END
  END PWDATA[5]
  PIN PWDATA[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 109.9500 21.5625 110.4600 21.6375 ;
    END
  END PWDATA[4]
  PIN PWDATA[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 109.9500 28.7625 110.4600 28.8375 ;
    END
  END PWDATA[3]
  PIN PWDATA[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 109.9500 22.4625 110.4600 22.5375 ;
    END
  END PWDATA[2]
  PIN PWDATA[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 109.9500 27.8625 110.4600 27.9375 ;
    END
  END PWDATA[1]
  PIN PWDATA[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 67.7625 0.0000 67.8375 0.5100 ;
    END
  END PWDATA[0]
  PIN PRDATA[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 109.9500 7.6125 110.4600 7.6875 ;
    END
  END PRDATA[31]
  PIN PRDATA[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 109.9500 7.3125 110.4600 7.3875 ;
    END
  END PRDATA[30]
  PIN PRDATA[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 109.9500 7.0125 110.4600 7.0875 ;
    END
  END PRDATA[29]
  PIN PRDATA[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 109.9500 6.7125 110.4600 6.7875 ;
    END
  END PRDATA[28]
  PIN PRDATA[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 109.9500 6.4125 110.4600 6.4875 ;
    END
  END PRDATA[27]
  PIN PRDATA[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 109.9500 6.1125 110.4600 6.1875 ;
    END
  END PRDATA[26]
  PIN PRDATA[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 109.9500 5.8125 110.4600 5.8875 ;
    END
  END PRDATA[25]
  PIN PRDATA[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 109.9500 5.5125 110.4600 5.5875 ;
    END
  END PRDATA[24]
  PIN PRDATA[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 109.9500 5.2125 110.4600 5.2875 ;
    END
  END PRDATA[23]
  PIN PRDATA[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 109.9500 4.9125 110.4600 4.9875 ;
    END
  END PRDATA[22]
  PIN PRDATA[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 109.9500 4.6125 110.4600 4.6875 ;
    END
  END PRDATA[21]
  PIN PRDATA[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 109.9500 4.3125 110.4600 4.3875 ;
    END
  END PRDATA[20]
  PIN PRDATA[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 109.9500 4.0125 110.4600 4.0875 ;
    END
  END PRDATA[19]
  PIN PRDATA[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 109.9500 3.7125 110.4600 3.7875 ;
    END
  END PRDATA[18]
  PIN PRDATA[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 109.9500 3.4125 110.4600 3.4875 ;
    END
  END PRDATA[17]
  PIN PRDATA[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 109.9500 3.1125 110.4600 3.1875 ;
    END
  END PRDATA[16]
  PIN PRDATA[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 109.9500 2.8125 110.4600 2.8875 ;
    END
  END PRDATA[15]
  PIN PRDATA[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 109.9500 2.5125 110.4600 2.5875 ;
    END
  END PRDATA[14]
  PIN PRDATA[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 109.9500 2.2125 110.4600 2.2875 ;
    END
  END PRDATA[13]
  PIN PRDATA[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 109.9500 1.9125 110.4600 1.9875 ;
    END
  END PRDATA[12]
  PIN PRDATA[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 109.9500 1.6125 110.4600 1.6875 ;
    END
  END PRDATA[11]
  PIN PRDATA[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 109.9500 1.3125 110.4600 1.3875 ;
    END
  END PRDATA[10]
  PIN PRDATA[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 109.9500 1.0125 110.4600 1.0875 ;
    END
  END PRDATA[9]
  PIN PRDATA[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 109.9500 1.0125 110.4600 1.0875 ;
    END
  END PRDATA[8]
  PIN PRDATA[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 67.2675 0.0000 67.3425 0.4200 ;
    END
  END PRDATA[7]
  PIN PRDATA[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 72.9375 0.0000 73.0125 0.4200 ;
    END
  END PRDATA[6]
  PIN PRDATA[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 70.8375 0.0000 70.9125 0.4200 ;
    END
  END PRDATA[5]
  PIN PRDATA[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 72.0975 0.0000 72.1725 0.4200 ;
    END
  END PRDATA[4]
  PIN PRDATA[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 65.3775 0.0000 65.4525 0.4200 ;
    END
  END PRDATA[3]
  PIN PRDATA[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 65.7975 0.0000 65.8725 0.4200 ;
    END
  END PRDATA[2]
  PIN PRDATA[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 67.6875 0.0000 67.7625 0.4200 ;
    END
  END PRDATA[1]
  PIN PRDATA[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 69.9975 0.0000 70.0725 0.4200 ;
    END
  END PRDATA[0]
  PIN PREADY
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 109.6125 0.0000 109.6875 0.5100 ;
    END
  END PREADY
  PIN PSLVERR
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 109.9500 1.3125 110.4600 1.3875 ;
    END
  END PSLVERR
  PIN INT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 63.2625 0.0000 63.3375 0.5100 ;
    END
  END INT
  PIN OUT1N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 78.3975 0.0000 78.4725 0.4200 ;
    END
  END OUT1N
  PIN OUT2N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 78.8175 0.0000 78.8925 0.4200 ;
    END
  END OUT2N
  PIN RTSN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 81.3375 0.0000 81.4125 0.4200 ;
    END
  END RTSN
  PIN DTRN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 77.5575 0.0000 77.6325 0.4200 ;
    END
  END DTRN
  PIN CTSN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 109.9500 10.9125 110.4600 10.9875 ;
    END
  END CTSN
  PIN DSRN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 109.9500 6.7125 110.4600 6.7875 ;
    END
  END DSRN
  PIN DCDN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 109.9500 8.8125 110.4600 8.8875 ;
    END
  END DCDN
  PIN RIN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 104.8575 0.0000 104.9325 0.4200 ;
    END
  END RIN
  PIN SIN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 81.7575 0.0000 81.8325 0.4200 ;
    END
  END SIN
  PIN SOUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 79.6575 0.0000 79.7325 0.4200 ;
    END
  END SOUT
  OBS
    LAYER M1 ;
        RECT 0.0000 0.0000 110.4600 110.2500 ;
    LAYER M2 ;
        RECT 0.0000 0.0000 110.4600 110.2500 ;
    LAYER M3 ;
        RECT 0.0000 0.0000 110.4600 110.2500 ;
    LAYER M4 ;
        RECT 0.0000 0.0000 110.4600 110.2500 ;
    LAYER M5 ;
        RECT 0.0000 0.0000 110.4600 110.2500 ;
    LAYER M6 ;
        RECT 0.0000 0.0000 110.4600 110.2500 ;
    LAYER M7 ;
        RECT 0.0000 0.0000 110.4600 110.2500 ;
    LAYER M8 ;
        RECT 0.0000 0.0000 110.4600 110.2500 ;
  END
END apb_uart


VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO axi_spi_slave_wrap
  CLASS BLOCK ;
    SIZE 54.8100 BY 53.5500 ;
  FOREIGN axi_spi_slave_wrap 0.000000 0.000000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 34.0875 0.0000 34.1625 0.4200 ;
    END
  END clk_i
  PIN rst_ni
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 35.3475 0.0000 35.4225 0.4200 ;
    END
  END rst_ni
  PIN test_mode
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8.4675 53.1300 8.5425 53.5500 ;
    END
  END test_mode
  PIN axi_master.aw_valid
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 38.3625 0.0000 38.4375 0.5100 ;
    END
  END axi_master.aw_valid
  PIN axi_master.aw_addr[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 27.8625 0.5100 27.9375 ;
    END
  END axi_master.aw_addr[31]
  PIN axi_master.aw_addr[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 25.0125 0.5100 25.0875 ;
    END
  END axi_master.aw_addr[30]
  PIN axi_master.aw_addr[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 24.4125 0.5100 24.4875 ;
    END
  END axi_master.aw_addr[29]
  PIN axi_master.aw_addr[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 21.5625 0.5100 21.6375 ;
    END
  END axi_master.aw_addr[28]
  PIN axi_master.aw_addr[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 20.3625 0.5100 20.4375 ;
    END
  END axi_master.aw_addr[27]
  PIN axi_master.aw_addr[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 21.1125 0.5100 21.1875 ;
    END
  END axi_master.aw_addr[26]
  PIN axi_master.aw_addr[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 19.7625 0.5100 19.8375 ;
    END
  END axi_master.aw_addr[25]
  PIN axi_master.aw_addr[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 13.6125 0.5100 13.6875 ;
    END
  END axi_master.aw_addr[24]
  PIN axi_master.aw_addr[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 12.4125 0.5100 12.4875 ;
    END
  END axi_master.aw_addr[23]
  PIN axi_master.aw_addr[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 7.0125 0.5100 7.0875 ;
    END
  END axi_master.aw_addr[22]
  PIN axi_master.aw_addr[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 7.7625 0.5100 7.8375 ;
    END
  END axi_master.aw_addr[21]
  PIN axi_master.aw_addr[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7.7625 0.0000 7.8375 0.5100 ;
    END
  END axi_master.aw_addr[20]
  PIN axi_master.aw_addr[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8.2125 0.0000 8.2875 0.5100 ;
    END
  END axi_master.aw_addr[19]
  PIN axi_master.aw_addr[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10.7625 0.0000 10.8375 0.5100 ;
    END
  END axi_master.aw_addr[18]
  PIN axi_master.aw_addr[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11.6625 0.0000 11.7375 0.5100 ;
    END
  END axi_master.aw_addr[17]
  PIN axi_master.aw_addr[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14.5125 0.0000 14.5875 0.5100 ;
    END
  END axi_master.aw_addr[16]
  PIN axi_master.aw_addr[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15.1125 0.0000 15.1875 0.5100 ;
    END
  END axi_master.aw_addr[15]
  PIN axi_master.aw_addr[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18.2625 0.0000 18.3375 0.5100 ;
    END
  END axi_master.aw_addr[14]
  PIN axi_master.aw_addr[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 19.1625 0.0000 19.2375 0.5100 ;
    END
  END axi_master.aw_addr[13]
  PIN axi_master.aw_addr[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 21.8625 0.0000 21.9375 0.5100 ;
    END
  END axi_master.aw_addr[12]
  PIN axi_master.aw_addr[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 22.4625 0.0000 22.5375 0.5100 ;
    END
  END axi_master.aw_addr[11]
  PIN axi_master.aw_addr[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 25.9125 0.0000 25.9875 0.5100 ;
    END
  END axi_master.aw_addr[10]
  PIN axi_master.aw_addr[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 26.6625 0.0000 26.7375 0.5100 ;
    END
  END axi_master.aw_addr[9]
  PIN axi_master.aw_addr[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 27.5625 0.0000 27.6375 0.5100 ;
    END
  END axi_master.aw_addr[8]
  PIN axi_master.aw_addr[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 28.4625 0.0000 28.5375 0.5100 ;
    END
  END axi_master.aw_addr[7]
  PIN axi_master.aw_addr[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 31.9125 0.0000 31.9875 0.5100 ;
    END
  END axi_master.aw_addr[6]
  PIN axi_master.aw_addr[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 30.7125 0.0000 30.7875 0.5100 ;
    END
  END axi_master.aw_addr[5]
  PIN axi_master.aw_addr[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 27.1125 0.0000 27.1875 0.5100 ;
    END
  END axi_master.aw_addr[4]
  PIN axi_master.aw_addr[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 26.3625 0.0000 26.4375 0.5100 ;
    END
  END axi_master.aw_addr[3]
  PIN axi_master.aw_addr[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 25.4625 0.0000 25.5375 0.5100 ;
    END
  END axi_master.aw_addr[2]
  PIN axi_master.aw_addr[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 54.3000 28.0125 54.8100 28.0875 ;
    END
  END axi_master.aw_addr[1]
  PIN axi_master.aw_addr[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 29.5125 53.0400 29.5875 53.5500 ;
    END
  END axi_master.aw_addr[0]
  PIN axi_master.aw_prot[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 54.3000 1.6125 54.8100 1.6875 ;
    END
  END axi_master.aw_prot[2]
  PIN axi_master.aw_prot[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 54.3000 1.3125 54.8100 1.3875 ;
    END
  END axi_master.aw_prot[1]
  PIN axi_master.aw_prot[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 54.3000 1.0125 54.8100 1.0875 ;
    END
  END axi_master.aw_prot[0]
  PIN axi_master.aw_region[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 54.3000 1.0125 54.8100 1.0875 ;
    END
  END axi_master.aw_region[3]
  PIN axi_master.aw_region[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 54.3000 1.3125 54.8100 1.3875 ;
    END
  END axi_master.aw_region[2]
  PIN axi_master.aw_region[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 54.3000 1.6125 54.8100 1.6875 ;
    END
  END axi_master.aw_region[1]
  PIN axi_master.aw_region[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 54.3000 1.9125 54.8100 1.9875 ;
    END
  END axi_master.aw_region[0]
  PIN axi_master.aw_len[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 54.3000 2.2125 54.8100 2.2875 ;
    END
  END axi_master.aw_len[7]
  PIN axi_master.aw_len[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 54.3000 2.5125 54.8100 2.5875 ;
    END
  END axi_master.aw_len[6]
  PIN axi_master.aw_len[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 54.3000 2.8125 54.8100 2.8875 ;
    END
  END axi_master.aw_len[5]
  PIN axi_master.aw_len[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 54.3000 3.1125 54.8100 3.1875 ;
    END
  END axi_master.aw_len[4]
  PIN axi_master.aw_len[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 54.3000 3.4125 54.8100 3.4875 ;
    END
  END axi_master.aw_len[3]
  PIN axi_master.aw_len[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 54.3000 3.7125 54.8100 3.7875 ;
    END
  END axi_master.aw_len[2]
  PIN axi_master.aw_len[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 54.3000 4.0125 54.8100 4.0875 ;
    END
  END axi_master.aw_len[1]
  PIN axi_master.aw_len[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 54.3000 4.3125 54.8100 4.3875 ;
    END
  END axi_master.aw_len[0]
  PIN axi_master.aw_size[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 54.3000 4.6125 54.8100 4.6875 ;
    END
  END axi_master.aw_size[2]
  PIN axi_master.aw_size[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 3.2625 0.5100 3.3375 ;
    END
  END axi_master.aw_size[1]
  PIN axi_master.aw_size[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 54.3000 4.9125 54.8100 4.9875 ;
    END
  END axi_master.aw_size[0]
  PIN axi_master.aw_burst[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 54.3000 5.2125 54.8100 5.2875 ;
    END
  END axi_master.aw_burst[1]
  PIN axi_master.aw_burst[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 54.3000 5.5125 54.8100 5.5875 ;
    END
  END axi_master.aw_burst[0]
  PIN axi_master.aw_lock
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 54.3000 5.8125 54.8100 5.8875 ;
    END
  END axi_master.aw_lock
  PIN axi_master.aw_cache[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 54.3000 6.1125 54.8100 6.1875 ;
    END
  END axi_master.aw_cache[3]
  PIN axi_master.aw_cache[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 54.3000 6.4125 54.8100 6.4875 ;
    END
  END axi_master.aw_cache[2]
  PIN axi_master.aw_cache[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 54.3000 6.7125 54.8100 6.7875 ;
    END
  END axi_master.aw_cache[1]
  PIN axi_master.aw_cache[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 54.3000 7.0125 54.8100 7.0875 ;
    END
  END axi_master.aw_cache[0]
  PIN axi_master.aw_qos[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 54.3000 7.3125 54.8100 7.3875 ;
    END
  END axi_master.aw_qos[3]
  PIN axi_master.aw_qos[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 54.3000 7.6125 54.8100 7.6875 ;
    END
  END axi_master.aw_qos[2]
  PIN axi_master.aw_qos[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 54.3000 7.9125 54.8100 7.9875 ;
    END
  END axi_master.aw_qos[1]
  PIN axi_master.aw_qos[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 54.3000 8.2125 54.8100 8.2875 ;
    END
  END axi_master.aw_qos[0]
  PIN axi_master.aw_id[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 54.3000 8.5125 54.8100 8.5875 ;
    END
  END axi_master.aw_id[1]
  PIN axi_master.aw_id[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 2.9625 0.5100 3.0375 ;
    END
  END axi_master.aw_id[0]
  PIN axi_master.aw_user[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 54.3000 8.8125 54.8100 8.8875 ;
    END
  END axi_master.aw_user[0]
  PIN axi_master.aw_ready
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 38.0775 0.0000 38.1525 0.4200 ;
    END
  END axi_master.aw_ready
  PIN axi_master.ar_valid
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 35.2125 0.0000 35.2875 0.5100 ;
    END
  END axi_master.ar_valid
  PIN axi_master.ar_addr[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 28.1625 0.5100 28.2375 ;
    END
  END axi_master.ar_addr[31]
  PIN axi_master.ar_addr[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 25.3125 0.5100 25.3875 ;
    END
  END axi_master.ar_addr[30]
  PIN axi_master.ar_addr[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 24.7125 0.5100 24.7875 ;
    END
  END axi_master.ar_addr[29]
  PIN axi_master.ar_addr[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 21.8625 0.5100 21.9375 ;
    END
  END axi_master.ar_addr[28]
  PIN axi_master.ar_addr[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 20.6625 0.5100 20.7375 ;
    END
  END axi_master.ar_addr[27]
  PIN axi_master.ar_addr[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 21.1125 0.5100 21.1875 ;
    END
  END axi_master.ar_addr[26]
  PIN axi_master.ar_addr[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 20.0625 0.5100 20.1375 ;
    END
  END axi_master.ar_addr[25]
  PIN axi_master.ar_addr[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 13.9125 0.5100 13.9875 ;
    END
  END axi_master.ar_addr[24]
  PIN axi_master.ar_addr[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 12.7125 0.5100 12.7875 ;
    END
  END axi_master.ar_addr[23]
  PIN axi_master.ar_addr[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 7.3125 0.5100 7.3875 ;
    END
  END axi_master.ar_addr[22]
  PIN axi_master.ar_addr[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 8.0625 0.5100 8.1375 ;
    END
  END axi_master.ar_addr[21]
  PIN axi_master.ar_addr[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7.8375 0.0000 7.9125 0.4200 ;
    END
  END axi_master.ar_addr[20]
  PIN axi_master.ar_addr[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8.2575 0.0000 8.3325 0.4200 ;
    END
  END axi_master.ar_addr[19]
  PIN axi_master.ar_addr[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10.7775 0.0000 10.8525 0.4200 ;
    END
  END axi_master.ar_addr[18]
  PIN axi_master.ar_addr[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11.6175 0.0000 11.6925 0.4200 ;
    END
  END axi_master.ar_addr[17]
  PIN axi_master.ar_addr[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14.5575 0.0000 14.6325 0.4200 ;
    END
  END axi_master.ar_addr[16]
  PIN axi_master.ar_addr[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15.1875 0.0000 15.2625 0.4200 ;
    END
  END axi_master.ar_addr[15]
  PIN axi_master.ar_addr[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18.3375 0.0000 18.4125 0.4200 ;
    END
  END axi_master.ar_addr[14]
  PIN axi_master.ar_addr[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 19.1775 0.0000 19.2525 0.4200 ;
    END
  END axi_master.ar_addr[13]
  PIN axi_master.ar_addr[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 21.9075 0.0000 21.9825 0.4200 ;
    END
  END axi_master.ar_addr[12]
  PIN axi_master.ar_addr[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 22.5375 0.0000 22.6125 0.4200 ;
    END
  END axi_master.ar_addr[11]
  PIN axi_master.ar_addr[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 25.8975 0.0000 25.9725 0.4200 ;
    END
  END axi_master.ar_addr[10]
  PIN axi_master.ar_addr[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 26.7375 0.0000 26.8125 0.4200 ;
    END
  END axi_master.ar_addr[9]
  PIN axi_master.ar_addr[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 27.5775 0.0000 27.6525 0.4200 ;
    END
  END axi_master.ar_addr[8]
  PIN axi_master.ar_addr[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 28.4175 0.0000 28.4925 0.4200 ;
    END
  END axi_master.ar_addr[7]
  PIN axi_master.ar_addr[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 31.9875 0.0000 32.0625 0.4200 ;
    END
  END axi_master.ar_addr[6]
  PIN axi_master.ar_addr[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 30.7275 0.0000 30.8025 0.4200 ;
    END
  END axi_master.ar_addr[5]
  PIN axi_master.ar_addr[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 27.1575 0.0000 27.2325 0.4200 ;
    END
  END axi_master.ar_addr[4]
  PIN axi_master.ar_addr[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 26.3175 0.0000 26.3925 0.4200 ;
    END
  END axi_master.ar_addr[3]
  PIN axi_master.ar_addr[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 25.4775 0.0000 25.5525 0.4200 ;
    END
  END axi_master.ar_addr[2]
  PIN axi_master.ar_addr[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 54.3000 28.3125 54.8100 28.3875 ;
    END
  END axi_master.ar_addr[1]
  PIN axi_master.ar_addr[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 29.4675 53.1300 29.5425 53.5500 ;
    END
  END axi_master.ar_addr[0]
  PIN axi_master.ar_prot[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 54.3000 9.1125 54.8100 9.1875 ;
    END
  END axi_master.ar_prot[2]
  PIN axi_master.ar_prot[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 54.3000 9.4125 54.8100 9.4875 ;
    END
  END axi_master.ar_prot[1]
  PIN axi_master.ar_prot[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 54.3000 9.7125 54.8100 9.7875 ;
    END
  END axi_master.ar_prot[0]
  PIN axi_master.ar_region[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 54.3000 10.0125 54.8100 10.0875 ;
    END
  END axi_master.ar_region[3]
  PIN axi_master.ar_region[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 54.3000 10.3125 54.8100 10.3875 ;
    END
  END axi_master.ar_region[2]
  PIN axi_master.ar_region[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 54.3000 10.6125 54.8100 10.6875 ;
    END
  END axi_master.ar_region[1]
  PIN axi_master.ar_region[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 54.3000 10.9125 54.8100 10.9875 ;
    END
  END axi_master.ar_region[0]
  PIN axi_master.ar_len[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 54.3000 11.2125 54.8100 11.2875 ;
    END
  END axi_master.ar_len[7]
  PIN axi_master.ar_len[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 54.3000 11.5125 54.8100 11.5875 ;
    END
  END axi_master.ar_len[6]
  PIN axi_master.ar_len[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 54.3000 11.8125 54.8100 11.8875 ;
    END
  END axi_master.ar_len[5]
  PIN axi_master.ar_len[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 54.3000 12.1125 54.8100 12.1875 ;
    END
  END axi_master.ar_len[4]
  PIN axi_master.ar_len[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 54.3000 12.4125 54.8100 12.4875 ;
    END
  END axi_master.ar_len[3]
  PIN axi_master.ar_len[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 54.3000 12.7125 54.8100 12.7875 ;
    END
  END axi_master.ar_len[2]
  PIN axi_master.ar_len[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 54.3000 13.0125 54.8100 13.0875 ;
    END
  END axi_master.ar_len[1]
  PIN axi_master.ar_len[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 54.3000 13.3125 54.8100 13.3875 ;
    END
  END axi_master.ar_len[0]
  PIN axi_master.ar_size[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 54.3000 13.6125 54.8100 13.6875 ;
    END
  END axi_master.ar_size[2]
  PIN axi_master.ar_size[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 2.6625 0.5100 2.7375 ;
    END
  END axi_master.ar_size[1]
  PIN axi_master.ar_size[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 54.3000 13.9125 54.8100 13.9875 ;
    END
  END axi_master.ar_size[0]
  PIN axi_master.ar_burst[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 54.3000 14.2125 54.8100 14.2875 ;
    END
  END axi_master.ar_burst[1]
  PIN axi_master.ar_burst[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 54.3000 14.5125 54.8100 14.5875 ;
    END
  END axi_master.ar_burst[0]
  PIN axi_master.ar_lock
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 54.3000 14.8125 54.8100 14.8875 ;
    END
  END axi_master.ar_lock
  PIN axi_master.ar_cache[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 54.3000 15.1125 54.8100 15.1875 ;
    END
  END axi_master.ar_cache[3]
  PIN axi_master.ar_cache[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 54.3000 15.4125 54.8100 15.4875 ;
    END
  END axi_master.ar_cache[2]
  PIN axi_master.ar_cache[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 54.3000 15.7125 54.8100 15.7875 ;
    END
  END axi_master.ar_cache[1]
  PIN axi_master.ar_cache[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 54.3000 16.0125 54.8100 16.0875 ;
    END
  END axi_master.ar_cache[0]
  PIN axi_master.ar_qos[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 54.3000 16.3125 54.8100 16.3875 ;
    END
  END axi_master.ar_qos[3]
  PIN axi_master.ar_qos[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 54.3000 16.6125 54.8100 16.6875 ;
    END
  END axi_master.ar_qos[2]
  PIN axi_master.ar_qos[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 54.3000 16.9125 54.8100 16.9875 ;
    END
  END axi_master.ar_qos[1]
  PIN axi_master.ar_qos[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 54.3000 17.2125 54.8100 17.2875 ;
    END
  END axi_master.ar_qos[0]
  PIN axi_master.ar_id[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 54.3000 17.5125 54.8100 17.5875 ;
    END
  END axi_master.ar_id[1]
  PIN axi_master.ar_id[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 2.3625 0.5100 2.4375 ;
    END
  END axi_master.ar_id[0]
  PIN axi_master.ar_user[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 54.3000 17.8125 54.8100 17.8875 ;
    END
  END axi_master.ar_user[0]
  PIN axi_master.ar_ready
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 35.5125 0.0000 35.5875 0.5100 ;
    END
  END axi_master.ar_ready
  PIN axi_master.w_valid
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 39.2625 0.0000 39.3375 0.5100 ;
    END
  END axi_master.w_valid
  PIN axi_master.w_data[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 54.3000 10.4625 54.8100 10.5375 ;
    END
  END axi_master.w_data[31]
  PIN axi_master.w_data[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 54.3000 8.3625 54.8100 8.4375 ;
    END
  END axi_master.w_data[30]
  PIN axi_master.w_data[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 54.3000 11.5125 54.8100 11.5875 ;
    END
  END axi_master.w_data[29]
  PIN axi_master.w_data[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 54.3000 12.5625 54.8100 12.6375 ;
    END
  END axi_master.w_data[28]
  PIN axi_master.w_data[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 47.3175 0.0000 47.3925 0.4200 ;
    END
  END axi_master.w_data[27]
  PIN axi_master.w_data[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 41.2275 0.0000 41.3025 0.4200 ;
    END
  END axi_master.w_data[26]
  PIN axi_master.w_data[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 54.3000 15.7125 54.8100 15.7875 ;
    END
  END axi_master.w_data[25]
  PIN axi_master.w_data[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 54.3000 6.2625 54.8100 6.3375 ;
    END
  END axi_master.w_data[24]
  PIN axi_master.w_data[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 41.8575 0.0000 41.9325 0.4200 ;
    END
  END axi_master.w_data[23]
  PIN axi_master.w_data[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 51.5175 0.0000 51.5925 0.4200 ;
    END
  END axi_master.w_data[22]
  PIN axi_master.w_data[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 54.3000 13.6125 54.8100 13.6875 ;
    END
  END axi_master.w_data[21]
  PIN axi_master.w_data[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 54.3000 13.3125 54.8100 13.3875 ;
    END
  END axi_master.w_data[20]
  PIN axi_master.w_data[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 54.3000 6.5625 54.8100 6.6375 ;
    END
  END axi_master.w_data[19]
  PIN axi_master.w_data[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 42.2775 0.0000 42.3525 0.4200 ;
    END
  END axi_master.w_data[18]
  PIN axi_master.w_data[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 54.3000 17.8125 54.8100 17.8875 ;
    END
  END axi_master.w_data[17]
  PIN axi_master.w_data[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 48.7875 0.0000 48.8625 0.4200 ;
    END
  END axi_master.w_data[16]
  PIN axi_master.w_data[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 54.3000 12.2625 54.8100 12.3375 ;
    END
  END axi_master.w_data[15]
  PIN axi_master.w_data[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 44.5875 0.0000 44.6625 0.4200 ;
    END
  END axi_master.w_data[14]
  PIN axi_master.w_data[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 44.6625 0.0000 44.7375 0.5100 ;
    END
  END axi_master.w_data[13]
  PIN axi_master.w_data[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 54.3000 9.4125 54.8100 9.4875 ;
    END
  END axi_master.w_data[12]
  PIN axi_master.w_data[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 46.6875 0.0000 46.7625 0.4200 ;
    END
  END axi_master.w_data[11]
  PIN axi_master.w_data[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 52.3575 0.0000 52.4325 0.4200 ;
    END
  END axi_master.w_data[10]
  PIN axi_master.w_data[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 45.0075 0.0000 45.0825 0.4200 ;
    END
  END axi_master.w_data[9]
  PIN axi_master.w_data[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 54.3000 11.2125 54.8100 11.2875 ;
    END
  END axi_master.w_data[8]
  PIN axi_master.w_data[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 54.3000 15.4125 54.8100 15.4875 ;
    END
  END axi_master.w_data[7]
  PIN axi_master.w_data[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 54.3000 4.1625 54.8100 4.2375 ;
    END
  END axi_master.w_data[6]
  PIN axi_master.w_data[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 45.4275 0.0000 45.5025 0.4200 ;
    END
  END axi_master.w_data[5]
  PIN axi_master.w_data[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 54.3000 8.0625 54.8100 8.1375 ;
    END
  END axi_master.w_data[4]
  PIN axi_master.w_data[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 54.3000 10.1625 54.8100 10.2375 ;
    END
  END axi_master.w_data[3]
  PIN axi_master.w_data[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 40.8075 0.0000 40.8825 0.4200 ;
    END
  END axi_master.w_data[2]
  PIN axi_master.w_data[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 48.7125 0.0000 48.7875 0.5100 ;
    END
  END axi_master.w_data[1]
  PIN axi_master.w_data[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 43.9575 0.0000 44.0325 0.4200 ;
    END
  END axi_master.w_data[0]
  PIN axi_master.w_strb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 2.0625 0.5100 2.1375 ;
    END
  END axi_master.w_strb[3]
  PIN axi_master.w_strb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1.7625 0.5100 1.8375 ;
    END
  END axi_master.w_strb[2]
  PIN axi_master.w_strb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1.4625 0.5100 1.5375 ;
    END
  END axi_master.w_strb[1]
  PIN axi_master.w_strb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1.1625 0.5100 1.2375 ;
    END
  END axi_master.w_strb[0]
  PIN axi_master.w_user[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 54.3000 18.1125 54.8100 18.1875 ;
    END
  END axi_master.w_user[0]
  PIN axi_master.w_last
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 0.8625 0.5100 0.9375 ;
    END
  END axi_master.w_last
  PIN axi_master.w_ready
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 38.9625 0.0000 39.0375 0.5100 ;
    END
  END axi_master.w_ready
  PIN axi_master.r_valid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 33.7125 0.0000 33.7875 0.5100 ;
    END
  END axi_master.r_valid
  PIN axi_master.r_data[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 34.5075 0.0000 34.5825 0.4200 ;
    END
  END axi_master.r_data[31]
  PIN axi_master.r_data[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 39.9675 0.0000 40.0425 0.4200 ;
    END
  END axi_master.r_data[30]
  PIN axi_master.r_data[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 37.6575 0.0000 37.7325 0.4200 ;
    END
  END axi_master.r_data[29]
  PIN axi_master.r_data[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 33.2475 0.0000 33.3225 0.4200 ;
    END
  END axi_master.r_data[28]
  PIN axi_master.r_data[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14.8125 0.0000 14.8875 0.5100 ;
    END
  END axi_master.r_data[27]
  PIN axi_master.r_data[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 32.6175 0.0000 32.6925 0.4200 ;
    END
  END axi_master.r_data[26]
  PIN axi_master.r_data[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 24.8475 0.0000 24.9225 0.4200 ;
    END
  END axi_master.r_data[25]
  PIN axi_master.r_data[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 23.7975 0.0000 23.8725 0.4200 ;
    END
  END axi_master.r_data[24]
  PIN axi_master.r_data[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 32.8125 0.0000 32.8875 0.5100 ;
    END
  END axi_master.r_data[23]
  PIN axi_master.r_data[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11.1975 0.0000 11.2725 0.4200 ;
    END
  END axi_master.r_data[22]
  PIN axi_master.r_data[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 30.3075 0.0000 30.3825 0.4200 ;
    END
  END axi_master.r_data[21]
  PIN axi_master.r_data[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17.9175 0.0000 17.9925 0.4200 ;
    END
  END axi_master.r_data[20]
  PIN axi_master.r_data[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 29.6775 0.0000 29.7525 0.4200 ;
    END
  END axi_master.r_data[19]
  PIN axi_master.r_data[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 38.9175 0.0000 38.9925 0.4200 ;
    END
  END axi_master.r_data[18]
  PIN axi_master.r_data[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 36.8175 0.0000 36.8925 0.4200 ;
    END
  END axi_master.r_data[17]
  PIN axi_master.r_data[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 39.5475 0.0000 39.6225 0.4200 ;
    END
  END axi_master.r_data[16]
  PIN axi_master.r_data[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15.6075 0.0000 15.6825 0.4200 ;
    END
  END axi_master.r_data[15]
  PIN axi_master.r_data[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 21.2775 0.0000 21.3525 0.4200 ;
    END
  END axi_master.r_data[14]
  PIN axi_master.r_data[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 36.1875 0.0000 36.2625 0.4200 ;
    END
  END axi_master.r_data[13]
  PIN axi_master.r_data[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 26.9625 0.0000 27.0375 0.5100 ;
    END
  END axi_master.r_data[12]
  PIN axi_master.r_data[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 35.7675 0.0000 35.8425 0.4200 ;
    END
  END axi_master.r_data[11]
  PIN axi_master.r_data[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18.7575 0.0000 18.8325 0.4200 ;
    END
  END axi_master.r_data[10]
  PIN axi_master.r_data[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 30.4125 0.0000 30.4875 0.5100 ;
    END
  END axi_master.r_data[9]
  PIN axi_master.r_data[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11.3625 0.0000 11.4375 0.5100 ;
    END
  END axi_master.r_data[8]
  PIN axi_master.r_data[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 33.6675 0.0000 33.7425 0.4200 ;
    END
  END axi_master.r_data[7]
  PIN axi_master.r_data[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 29.2575 0.0000 29.3325 0.4200 ;
    END
  END axi_master.r_data[6]
  PIN axi_master.r_data[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 26.0625 0.0000 26.1375 0.5100 ;
    END
  END axi_master.r_data[5]
  PIN axi_master.r_data[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 22.9575 0.0000 23.0325 0.4200 ;
    END
  END axi_master.r_data[4]
  PIN axi_master.r_data[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 21.2625 0.0000 21.3375 0.5100 ;
    END
  END axi_master.r_data[3]
  PIN axi_master.r_data[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 26.6625 0.0000 26.7375 0.5100 ;
    END
  END axi_master.r_data[2]
  PIN axi_master.r_data[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 40.3875 0.0000 40.4625 0.4200 ;
    END
  END axi_master.r_data[1]
  PIN axi_master.r_data[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 27.9975 0.0000 28.0725 0.4200 ;
    END
  END axi_master.r_data[0]
  PIN axi_master.r_resp[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 27.7125 53.0400 27.7875 53.5500 ;
    END
  END axi_master.r_resp[1]
  PIN axi_master.r_resp[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 27.7125 53.0400 27.7875 53.5500 ;
    END
  END axi_master.r_resp[0]
  PIN axi_master.r_last
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 26.9475 53.1300 27.0225 53.5500 ;
    END
  END axi_master.r_last
  PIN axi_master.r_id[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 27.1125 53.0400 27.1875 53.5500 ;
    END
  END axi_master.r_id[1]
  PIN axi_master.r_id[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 27.7875 53.1300 27.8625 53.5500 ;
    END
  END axi_master.r_id[0]
  PIN axi_master.r_user[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 27.7125 0.0000 27.7875 0.5100 ;
    END
  END axi_master.r_user[0]
  PIN axi_master.r_ready
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 33.4125 0.0000 33.4875 0.5100 ;
    END
  END axi_master.r_ready
  PIN axi_master.b_valid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 40.6125 0.0000 40.6875 0.5100 ;
    END
  END axi_master.b_valid
  PIN axi_master.b_resp[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 27.4125 53.0400 27.4875 53.5500 ;
    END
  END axi_master.b_resp[1]
  PIN axi_master.b_resp[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 27.4125 0.0000 27.4875 0.5100 ;
    END
  END axi_master.b_resp[0]
  PIN axi_master.b_id[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 27.3675 53.1300 27.4425 53.5500 ;
    END
  END axi_master.b_id[1]
  PIN axi_master.b_id[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 27.4125 53.0400 27.4875 53.5500 ;
    END
  END axi_master.b_id[0]
  PIN axi_master.b_user[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 27.1125 53.0400 27.1875 53.5500 ;
    END
  END axi_master.b_user[0]
  PIN axi_master.b_ready
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 41.3625 0.0000 41.4375 0.5100 ;
    END
  END axi_master.b_ready
  PIN spi_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 23.3775 53.1300 23.4525 53.5500 ;
    END
  END spi_clk
  PIN spi_cs
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 28.8375 0.0000 28.9125 0.4200 ;
    END
  END spi_cs
  PIN spi_mode[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 33.0375 53.1300 33.1125 53.5500 ;
    END
  END spi_mode[1]
  PIN spi_mode[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 35.1375 53.1300 35.2125 53.5500 ;
    END
  END spi_mode[0]
  PIN spi_sdo0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15.3975 53.1300 15.4725 53.5500 ;
    END
  END spi_sdo0
  PIN spi_sdo1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13.5075 53.1300 13.5825 53.5500 ;
    END
  END spi_sdo1
  PIN spi_sdo2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14.1375 53.1300 14.2125 53.5500 ;
    END
  END spi_sdo2
  PIN spi_sdo3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15.5625 53.0400 15.6375 53.5500 ;
    END
  END spi_sdo3
  PIN spi_sdi0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 28.0125 0.5100 28.0875 ;
    END
  END spi_sdi0
  PIN spi_sdi1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 28.9125 0.5100 28.9875 ;
    END
  END spi_sdi1
  PIN spi_sdi2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 28.6125 0.5100 28.6875 ;
    END
  END spi_sdi2
  PIN spi_sdi3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 25.6125 0.5100 25.6875 ;
    END
  END spi_sdi3
  OBS
    LAYER M1 ;
        RECT 0.0000 0.0000 54.8100 53.5500 ;
    LAYER M2 ;
        RECT 0.0000 0.0000 54.8100 53.5500 ;
    LAYER M3 ;
        RECT 0.0000 0.0000 54.8100 53.5500 ;
    LAYER M4 ;
        RECT 0.0000 0.0000 54.8100 53.5500 ;
    LAYER M5 ;
        RECT 0.0000 0.0000 54.8100 53.5500 ;
    LAYER M6 ;
        RECT 0.0000 0.0000 54.8100 53.5500 ;
    LAYER M7 ;
        RECT 0.0000 0.0000 54.8100 53.5500 ;
    LAYER M8 ;
        RECT 0.0000 0.0000 54.8100 53.5500 ;
  END
END axi_spi_slave_wrap


VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO periph_bus_wrap
  CLASS BLOCK ;
    SIZE 40.3200 BY 39.9000 ;
  FOREIGN periph_bus_wrap 0.000000 0.000000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 20.0175 39.4800 20.0925 39.9000 ;
    END
  END clk_i
  PIN rst_ni
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 21.7125 0.0000 21.7875 0.5100 ;
    END
  END rst_ni
  PIN apb_slave.paddr[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 4.6125 0.5100 4.6875 ;
    END
  END apb_slave.paddr[31]
  PIN apb_slave.paddr[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9.9375 0.0000 10.0125 0.4200 ;
    END
  END apb_slave.paddr[30]
  PIN apb_slave.paddr[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8.8875 0.0000 8.9625 0.4200 ;
    END
  END apb_slave.paddr[29]
  PIN apb_slave.paddr[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13.7175 0.0000 13.7925 0.4200 ;
    END
  END apb_slave.paddr[28]
  PIN apb_slave.paddr[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16.0275 0.0000 16.1025 0.4200 ;
    END
  END apb_slave.paddr[27]
  PIN apb_slave.paddr[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 5.6625 0.5100 5.7375 ;
    END
  END apb_slave.paddr[26]
  PIN apb_slave.paddr[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16.1625 0.0000 16.2375 0.5100 ;
    END
  END apb_slave.paddr[25]
  PIN apb_slave.paddr[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7.8375 0.0000 7.9125 0.4200 ;
    END
  END apb_slave.paddr[24]
  PIN apb_slave.paddr[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 3.1125 0.5100 3.1875 ;
    END
  END apb_slave.paddr[23]
  PIN apb_slave.paddr[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7.9125 0.0000 7.9875 0.5100 ;
    END
  END apb_slave.paddr[22]
  PIN apb_slave.paddr[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10.9875 0.0000 11.0625 0.4200 ;
    END
  END apb_slave.paddr[21]
  PIN apb_slave.paddr[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17.2875 0.0000 17.3625 0.4200 ;
    END
  END apb_slave.paddr[20]
  PIN apb_slave.paddr[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 25.2675 0.0000 25.3425 0.4200 ;
    END
  END apb_slave.paddr[19]
  PIN apb_slave.paddr[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.8100 5.8125 40.3200 5.8875 ;
    END
  END apb_slave.paddr[18]
  PIN apb_slave.paddr[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 29.2575 0.0000 29.3325 0.4200 ;
    END
  END apb_slave.paddr[17]
  PIN apb_slave.paddr[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 33.8775 0.0000 33.9525 0.4200 ;
    END
  END apb_slave.paddr[16]
  PIN apb_slave.paddr[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 30.9375 0.0000 31.0125 0.4200 ;
    END
  END apb_slave.paddr[15]
  PIN apb_slave.paddr[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 27.3675 0.0000 27.4425 0.4200 ;
    END
  END apb_slave.paddr[14]
  PIN apb_slave.paddr[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 24.2175 0.0000 24.2925 0.4200 ;
    END
  END apb_slave.paddr[13]
  PIN apb_slave.paddr[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 24.7125 0.0000 24.7875 0.5100 ;
    END
  END apb_slave.paddr[12]
  PIN apb_slave.paddr[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8.0475 39.4800 8.1225 39.9000 ;
    END
  END apb_slave.paddr[11]
  PIN apb_slave.paddr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 22.6125 0.5100 22.6875 ;
    END
  END apb_slave.paddr[10]
  PIN apb_slave.paddr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9.5175 39.4800 9.5925 39.9000 ;
    END
  END apb_slave.paddr[9]
  PIN apb_slave.paddr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14.1375 39.4800 14.2125 39.9000 ;
    END
  END apb_slave.paddr[8]
  PIN apb_slave.paddr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 27.5625 0.5100 27.6375 ;
    END
  END apb_slave.paddr[7]
  PIN apb_slave.paddr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14.5575 39.4800 14.6325 39.9000 ;
    END
  END apb_slave.paddr[6]
  PIN apb_slave.paddr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 22.3125 0.5100 22.3875 ;
    END
  END apb_slave.paddr[5]
  PIN apb_slave.paddr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 12.7125 0.5100 12.7875 ;
    END
  END apb_slave.paddr[4]
  PIN apb_slave.paddr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 29.3625 0.5100 29.4375 ;
    END
  END apb_slave.paddr[3]
  PIN apb_slave.paddr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14.8125 39.3900 14.8875 39.9000 ;
    END
  END apb_slave.paddr[2]
  PIN apb_slave.paddr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12.0375 39.4800 12.1125 39.9000 ;
    END
  END apb_slave.paddr[1]
  PIN apb_slave.paddr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10.1475 39.4800 10.2225 39.9000 ;
    END
  END apb_slave.paddr[0]
  PIN apb_slave.pwdata[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 19.9125 0.5100 19.9875 ;
    END
  END apb_slave.pwdata[31]
  PIN apb_slave.pwdata[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 12.8625 0.5100 12.9375 ;
    END
  END apb_slave.pwdata[30]
  PIN apb_slave.pwdata[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 32.8125 0.5100 32.8875 ;
    END
  END apb_slave.pwdata[29]
  PIN apb_slave.pwdata[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 12.5625 0.5100 12.6375 ;
    END
  END apb_slave.pwdata[28]
  PIN apb_slave.pwdata[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18.3375 39.4800 18.4125 39.9000 ;
    END
  END apb_slave.pwdata[27]
  PIN apb_slave.pwdata[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 30.1125 0.5100 30.1875 ;
    END
  END apb_slave.pwdata[26]
  PIN apb_slave.pwdata[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12.2625 39.3900 12.3375 39.9000 ;
    END
  END apb_slave.pwdata[25]
  PIN apb_slave.pwdata[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 20.0625 39.3900 20.1375 39.9000 ;
    END
  END apb_slave.pwdata[24]
  PIN apb_slave.pwdata[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 23.3625 0.5100 23.4375 ;
    END
  END apb_slave.pwdata[23]
  PIN apb_slave.pwdata[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 27.4125 0.5100 27.4875 ;
    END
  END apb_slave.pwdata[22]
  PIN apb_slave.pwdata[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 25.1625 0.5100 25.2375 ;
    END
  END apb_slave.pwdata[21]
  PIN apb_slave.pwdata[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 21.8625 0.5100 21.9375 ;
    END
  END apb_slave.pwdata[20]
  PIN apb_slave.pwdata[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 20.3625 0.5100 20.4375 ;
    END
  END apb_slave.pwdata[19]
  PIN apb_slave.pwdata[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4.2675 39.4800 4.3425 39.9000 ;
    END
  END apb_slave.pwdata[18]
  PIN apb_slave.pwdata[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 19.9125 0.5100 19.9875 ;
    END
  END apb_slave.pwdata[17]
  PIN apb_slave.pwdata[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6.3675 39.4800 6.4425 39.9000 ;
    END
  END apb_slave.pwdata[16]
  PIN apb_slave.pwdata[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 22.4625 0.5100 22.5375 ;
    END
  END apb_slave.pwdata[15]
  PIN apb_slave.pwdata[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 19.3125 0.5100 19.3875 ;
    END
  END apb_slave.pwdata[14]
  PIN apb_slave.pwdata[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 17.0625 0.5100 17.1375 ;
    END
  END apb_slave.pwdata[13]
  PIN apb_slave.pwdata[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 20.9625 0.5100 21.0375 ;
    END
  END apb_slave.pwdata[12]
  PIN apb_slave.pwdata[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 22.9125 0.5100 22.9875 ;
    END
  END apb_slave.pwdata[11]
  PIN apb_slave.pwdata[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 12.4125 0.5100 12.4875 ;
    END
  END apb_slave.pwdata[10]
  PIN apb_slave.pwdata[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 27.2625 0.5100 27.3375 ;
    END
  END apb_slave.pwdata[9]
  PIN apb_slave.pwdata[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16.4475 39.4800 16.5225 39.9000 ;
    END
  END apb_slave.pwdata[8]
  PIN apb_slave.pwdata[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 18.2625 0.5100 18.3375 ;
    END
  END apb_slave.pwdata[7]
  PIN apb_slave.pwdata[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 13.9125 0.0000 13.9875 0.5100 ;
    END
  END apb_slave.pwdata[6]
  PIN apb_slave.pwdata[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 19.5975 39.4800 19.6725 39.9000 ;
    END
  END apb_slave.pwdata[5]
  PIN apb_slave.pwdata[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 12.2625 0.5100 12.3375 ;
    END
  END apb_slave.pwdata[4]
  PIN apb_slave.pwdata[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 12.1125 0.5100 12.1875 ;
    END
  END apb_slave.pwdata[3]
  PIN apb_slave.pwdata[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 17.6625 0.5100 17.7375 ;
    END
  END apb_slave.pwdata[2]
  PIN apb_slave.pwdata[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 13.0125 0.5100 13.0875 ;
    END
  END apb_slave.pwdata[1]
  PIN apb_slave.pwdata[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 27.1125 0.5100 27.1875 ;
    END
  END apb_slave.pwdata[0]
  PIN apb_slave.pwrite
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 4.3125 0.5100 4.3875 ;
    END
  END apb_slave.pwrite
  PIN apb_slave.psel
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 21.8625 0.0000 21.9375 0.5100 ;
    END
  END apb_slave.psel
  PIN apb_slave.penable
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 4.0125 0.5100 4.0875 ;
    END
  END apb_slave.penable
  PIN apb_slave.prdata[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 21.2625 39.3900 21.3375 39.9000 ;
    END
  END apb_slave.prdata[31]
  PIN apb_slave.prdata[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 24.2175 39.4800 24.2925 39.9000 ;
    END
  END apb_slave.prdata[30]
  PIN apb_slave.prdata[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.8100 31.1625 40.3200 31.2375 ;
    END
  END apb_slave.prdata[29]
  PIN apb_slave.prdata[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.8100 19.1625 40.3200 19.2375 ;
    END
  END apb_slave.prdata[28]
  PIN apb_slave.prdata[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 38.1975 12.9000 40.3200 13.5000 ;
    END
  END apb_slave.prdata[27]
  PIN apb_slave.prdata[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 22.7475 39.4800 22.8225 39.9000 ;
    END
  END apb_slave.prdata[26]
  PIN apb_slave.prdata[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 27.7875 39.4800 27.8625 39.9000 ;
    END
  END apb_slave.prdata[25]
  PIN apb_slave.prdata[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.8100 25.4625 40.3200 25.5375 ;
    END
  END apb_slave.prdata[24]
  PIN apb_slave.prdata[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.8100 25.1625 40.3200 25.2375 ;
    END
  END apb_slave.prdata[23]
  PIN apb_slave.prdata[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.8100 27.5625 40.3200 27.6375 ;
    END
  END apb_slave.prdata[22]
  PIN apb_slave.prdata[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.8100 17.0625 40.3200 17.1375 ;
    END
  END apb_slave.prdata[21]
  PIN apb_slave.prdata[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.8100 29.0625 40.3200 29.1375 ;
    END
  END apb_slave.prdata[20]
  PIN apb_slave.prdata[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.8100 33.2625 40.3200 33.3375 ;
    END
  END apb_slave.prdata[19]
  PIN apb_slave.prdata[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.8100 22.7625 40.3200 22.8375 ;
    END
  END apb_slave.prdata[18]
  PIN apb_slave.prdata[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.8100 21.2625 40.3200 21.3375 ;
    END
  END apb_slave.prdata[17]
  PIN apb_slave.prdata[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 24.6375 39.4800 24.7125 39.9000 ;
    END
  END apb_slave.prdata[16]
  PIN apb_slave.prdata[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 38.1975 18.9000 40.3200 19.5000 ;
    END
  END apb_slave.prdata[15]
  PIN apb_slave.prdata[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 21.0675 0.0000 21.1425 0.4200 ;
    END
  END apb_slave.prdata[14]
  PIN apb_slave.prdata[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.8100 11.5125 40.3200 11.5875 ;
    END
  END apb_slave.prdata[13]
  PIN apb_slave.prdata[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 32.1975 39.4800 32.2725 39.9000 ;
    END
  END apb_slave.prdata[12]
  PIN apb_slave.prdata[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 38.1975 22.5000 40.3200 23.1000 ;
    END
  END apb_slave.prdata[11]
  PIN apb_slave.prdata[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 20.2125 39.3900 20.2875 39.9000 ;
    END
  END apb_slave.prdata[10]
  PIN apb_slave.prdata[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.8100 20.6625 40.3200 20.7375 ;
    END
  END apb_slave.prdata[9]
  PIN apb_slave.prdata[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 16.9125 39.3900 16.9875 39.9000 ;
    END
  END apb_slave.prdata[8]
  PIN apb_slave.prdata[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 36.1875 39.4800 36.2625 39.9000 ;
    END
  END apb_slave.prdata[7]
  PIN apb_slave.prdata[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.8100 24.8625 40.3200 24.9375 ;
    END
  END apb_slave.prdata[6]
  PIN apb_slave.prdata[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 21.7125 39.3900 21.7875 39.9000 ;
    END
  END apb_slave.prdata[5]
  PIN apb_slave.prdata[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 25.8975 39.4800 25.9725 39.9000 ;
    END
  END apb_slave.prdata[4]
  PIN apb_slave.prdata[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.8100 25.7625 40.3200 25.8375 ;
    END
  END apb_slave.prdata[3]
  PIN apb_slave.prdata[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 33.4575 39.4800 33.5325 39.9000 ;
    END
  END apb_slave.prdata[2]
  PIN apb_slave.prdata[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 29.8875 39.4800 29.9625 39.9000 ;
    END
  END apb_slave.prdata[1]
  PIN apb_slave.prdata[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.8100 14.9625 40.3200 15.0375 ;
    END
  END apb_slave.prdata[0]
  PIN apb_slave.pready
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 37.7625 0.0000 37.8375 0.5100 ;
    END
  END apb_slave.pready
  PIN apb_slave.pslverr
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 30.1125 0.0000 30.1875 0.5100 ;
    END
  END apb_slave.pslverr
  PIN uart_master.paddr[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 0.8625 40.3200 0.9375 ;
    END
  END uart_master.paddr[31]
  PIN uart_master.paddr[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 1.1625 40.3200 1.2375 ;
    END
  END uart_master.paddr[30]
  PIN uart_master.paddr[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 1.4625 40.3200 1.5375 ;
    END
  END uart_master.paddr[29]
  PIN uart_master.paddr[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 27.5625 0.0000 27.6375 0.5100 ;
    END
  END uart_master.paddr[28]
  PIN uart_master.paddr[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 27.8625 0.0000 27.9375 0.5100 ;
    END
  END uart_master.paddr[27]
  PIN uart_master.paddr[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 1.7625 40.3200 1.8375 ;
    END
  END uart_master.paddr[26]
  PIN uart_master.paddr[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 28.1625 0.0000 28.2375 0.5100 ;
    END
  END uart_master.paddr[25]
  PIN uart_master.paddr[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 2.0625 40.3200 2.1375 ;
    END
  END uart_master.paddr[24]
  PIN uart_master.paddr[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 2.3625 40.3200 2.4375 ;
    END
  END uart_master.paddr[23]
  PIN uart_master.paddr[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 2.6625 40.3200 2.7375 ;
    END
  END uart_master.paddr[22]
  PIN uart_master.paddr[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 2.9625 40.3200 3.0375 ;
    END
  END uart_master.paddr[21]
  PIN uart_master.paddr[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 28.4625 0.0000 28.5375 0.5100 ;
    END
  END uart_master.paddr[20]
  PIN uart_master.paddr[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 3.2625 40.3200 3.3375 ;
    END
  END uart_master.paddr[19]
  PIN uart_master.paddr[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 3.5625 40.3200 3.6375 ;
    END
  END uart_master.paddr[18]
  PIN uart_master.paddr[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 3.8625 40.3200 3.9375 ;
    END
  END uart_master.paddr[17]
  PIN uart_master.paddr[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 4.1625 40.3200 4.2375 ;
    END
  END uart_master.paddr[16]
  PIN uart_master.paddr[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 4.4625 40.3200 4.5375 ;
    END
  END uart_master.paddr[15]
  PIN uart_master.paddr[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 4.7625 40.3200 4.8375 ;
    END
  END uart_master.paddr[14]
  PIN uart_master.paddr[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 5.0625 40.3200 5.1375 ;
    END
  END uart_master.paddr[13]
  PIN uart_master.paddr[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 5.3625 40.3200 5.4375 ;
    END
  END uart_master.paddr[12]
  PIN uart_master.paddr[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1.9575 39.4800 2.0325 39.9000 ;
    END
  END uart_master.paddr[11]
  PIN uart_master.paddr[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7.4175 0.0000 7.4925 0.4200 ;
    END
  END uart_master.paddr[10]
  PIN uart_master.paddr[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 37.9125 0.5100 37.9875 ;
    END
  END uart_master.paddr[9]
  PIN uart_master.paddr[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 37.9125 0.5100 37.9875 ;
    END
  END uart_master.paddr[8]
  PIN uart_master.paddr[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1.9125 39.3900 1.9875 39.9000 ;
    END
  END uart_master.paddr[7]
  PIN uart_master.paddr[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 1.7625 39.3900 1.8375 39.9000 ;
    END
  END uart_master.paddr[6]
  PIN uart_master.paddr[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 9.8625 0.0000 9.9375 0.5100 ;
    END
  END uart_master.paddr[5]
  PIN uart_master.paddr[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7.4625 0.0000 7.5375 0.5100 ;
    END
  END uart_master.paddr[4]
  PIN uart_master.paddr[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 38.2125 0.5100 38.2875 ;
    END
  END uart_master.paddr[3]
  PIN uart_master.paddr[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 38.2125 0.5100 38.2875 ;
    END
  END uart_master.paddr[2]
  PIN uart_master.paddr[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1.5375 39.4800 1.6125 39.9000 ;
    END
  END uart_master.paddr[1]
  PIN uart_master.paddr[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1.6125 39.3900 1.6875 39.9000 ;
    END
  END uart_master.paddr[0]
  PIN uart_master.pwdata[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13.1625 0.0000 13.2375 0.5100 ;
    END
  END uart_master.pwdata[31]
  PIN uart_master.pwdata[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12.2475 0.0000 12.3225 0.4200 ;
    END
  END uart_master.pwdata[30]
  PIN uart_master.pwdata[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 38.8125 0.5100 38.8875 ;
    END
  END uart_master.pwdata[29]
  PIN uart_master.pwdata[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6.5775 0.0000 6.6525 0.4200 ;
    END
  END uart_master.pwdata[28]
  PIN uart_master.pwdata[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 38.8125 0.5100 38.8875 ;
    END
  END uart_master.pwdata[27]
  PIN uart_master.pwdata[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1.0125 39.3900 1.0875 39.9000 ;
    END
  END uart_master.pwdata[26]
  PIN uart_master.pwdata[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 0.8625 39.3900 0.9375 39.9000 ;
    END
  END uart_master.pwdata[25]
  PIN uart_master.pwdata[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 20.6625 0.0000 20.7375 0.5100 ;
    END
  END uart_master.pwdata[24]
  PIN uart_master.pwdata[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 5.5125 0.5100 5.5875 ;
    END
  END uart_master.pwdata[23]
  PIN uart_master.pwdata[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 10.6125 0.0000 10.6875 0.5100 ;
    END
  END uart_master.pwdata[22]
  PIN uart_master.pwdata[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 5.3625 0.5100 5.4375 ;
    END
  END uart_master.pwdata[21]
  PIN uart_master.pwdata[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 5.2125 0.5100 5.2875 ;
    END
  END uart_master.pwdata[20]
  PIN uart_master.pwdata[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 16.4625 0.0000 16.5375 0.5100 ;
    END
  END uart_master.pwdata[19]
  PIN uart_master.pwdata[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 5.0625 0.5100 5.1375 ;
    END
  END uart_master.pwdata[18]
  PIN uart_master.pwdata[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5.1075 0.0000 5.1825 0.4200 ;
    END
  END uart_master.pwdata[17]
  PIN uart_master.pwdata[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6.5625 0.0000 6.6375 0.5100 ;
    END
  END uart_master.pwdata[16]
  PIN uart_master.pwdata[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15.8625 0.0000 15.9375 0.5100 ;
    END
  END uart_master.pwdata[15]
  PIN uart_master.pwdata[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9.5625 0.0000 9.6375 0.5100 ;
    END
  END uart_master.pwdata[14]
  PIN uart_master.pwdata[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 15.7125 0.0000 15.7875 0.5100 ;
    END
  END uart_master.pwdata[13]
  PIN uart_master.pwdata[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7.1625 0.0000 7.2375 0.5100 ;
    END
  END uart_master.pwdata[12]
  PIN uart_master.pwdata[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12.1125 0.0000 12.1875 0.5100 ;
    END
  END uart_master.pwdata[11]
  PIN uart_master.pwdata[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 4.9125 0.5100 4.9875 ;
    END
  END uart_master.pwdata[10]
  PIN uart_master.pwdata[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5.0625 0.0000 5.1375 0.5100 ;
    END
  END uart_master.pwdata[9]
  PIN uart_master.pwdata[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 12.1125 0.0000 12.1875 0.5100 ;
    END
  END uart_master.pwdata[8]
  PIN uart_master.pwdata[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 8.6625 0.0000 8.7375 0.5100 ;
    END
  END uart_master.pwdata[7]
  PIN uart_master.pwdata[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11.8125 0.0000 11.8875 0.5100 ;
    END
  END uart_master.pwdata[6]
  PIN uart_master.pwdata[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 21.4125 0.0000 21.4875 0.5100 ;
    END
  END uart_master.pwdata[5]
  PIN uart_master.pwdata[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 9.2625 0.0000 9.3375 0.5100 ;
    END
  END uart_master.pwdata[4]
  PIN uart_master.pwdata[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 4.6125 0.5100 4.6875 ;
    END
  END uart_master.pwdata[3]
  PIN uart_master.pwdata[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5.3625 0.0000 5.4375 0.5100 ;
    END
  END uart_master.pwdata[2]
  PIN uart_master.pwdata[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 4.3125 0.5100 4.3875 ;
    END
  END uart_master.pwdata[1]
  PIN uart_master.pwdata[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 11.8125 0.0000 11.8875 0.5100 ;
    END
  END uart_master.pwdata[0]
  PIN uart_master.pwrite
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5.5275 0.0000 5.6025 0.4200 ;
    END
  END uart_master.pwrite
  PIN uart_master.psel
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 28.4175 0.0000 28.4925 0.4200 ;
    END
  END uart_master.psel
  PIN uart_master.penable
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 4.0125 0.5100 4.0875 ;
    END
  END uart_master.penable
  PIN uart_master.prdata[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 38.0625 39.3900 38.1375 39.9000 ;
    END
  END uart_master.prdata[31]
  PIN uart_master.prdata[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 37.7625 39.3900 37.8375 39.9000 ;
    END
  END uart_master.prdata[30]
  PIN uart_master.prdata[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 39.1125 39.3900 39.1875 39.9000 ;
    END
  END uart_master.prdata[29]
  PIN uart_master.prdata[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 37.4475 0.0000 37.5225 0.4200 ;
    END
  END uart_master.prdata[28]
  PIN uart_master.prdata[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 35.5125 0.0000 35.5875 0.5100 ;
    END
  END uart_master.prdata[27]
  PIN uart_master.prdata[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 38.3625 39.3900 38.4375 39.9000 ;
    END
  END uart_master.prdata[26]
  PIN uart_master.prdata[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 38.0625 39.3900 38.1375 39.9000 ;
    END
  END uart_master.prdata[25]
  PIN uart_master.prdata[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 38.3625 39.3900 38.4375 39.9000 ;
    END
  END uart_master.prdata[24]
  PIN uart_master.prdata[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 38.6625 39.3900 38.7375 39.9000 ;
    END
  END uart_master.prdata[23]
  PIN uart_master.prdata[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 38.8125 39.3900 38.8875 39.9000 ;
    END
  END uart_master.prdata[22]
  PIN uart_master.prdata[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 36.1125 0.0000 36.1875 0.5100 ;
    END
  END uart_master.prdata[21]
  PIN uart_master.prdata[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.8100 2.5125 40.3200 2.5875 ;
    END
  END uart_master.prdata[20]
  PIN uart_master.prdata[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.8100 2.2125 40.3200 2.2875 ;
    END
  END uart_master.prdata[19]
  PIN uart_master.prdata[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 37.0125 0.0000 37.0875 0.5100 ;
    END
  END uart_master.prdata[18]
  PIN uart_master.prdata[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 26.3625 0.0000 26.4375 0.5100 ;
    END
  END uart_master.prdata[17]
  PIN uart_master.prdata[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 26.0625 0.0000 26.1375 0.5100 ;
    END
  END uart_master.prdata[16]
  PIN uart_master.prdata[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 25.0125 0.0000 25.0875 0.5100 ;
    END
  END uart_master.prdata[15]
  PIN uart_master.prdata[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 21.9075 0.0000 21.9825 0.4200 ;
    END
  END uart_master.prdata[14]
  PIN uart_master.prdata[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 37.3125 0.0000 37.3875 0.5100 ;
    END
  END uart_master.prdata[13]
  PIN uart_master.prdata[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 1.4625 39.3900 1.5375 39.9000 ;
    END
  END uart_master.prdata[12]
  PIN uart_master.prdata[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 31.9875 0.0000 32.0625 0.4200 ;
    END
  END uart_master.prdata[11]
  PIN uart_master.prdata[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 38.5125 0.5100 38.5875 ;
    END
  END uart_master.prdata[10]
  PIN uart_master.prdata[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 37.4625 0.0000 37.5375 0.5100 ;
    END
  END uart_master.prdata[9]
  PIN uart_master.prdata[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 38.5125 0.5100 38.5875 ;
    END
  END uart_master.prdata[8]
  PIN uart_master.prdata[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 35.1375 0.0000 35.2125 0.4200 ;
    END
  END uart_master.prdata[7]
  PIN uart_master.prdata[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 36.7125 0.0000 36.7875 0.5100 ;
    END
  END uart_master.prdata[6]
  PIN uart_master.prdata[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 20.3625 0.0000 20.4375 0.5100 ;
    END
  END uart_master.prdata[5]
  PIN uart_master.prdata[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1.3125 39.3900 1.3875 39.9000 ;
    END
  END uart_master.prdata[4]
  PIN uart_master.prdata[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 37.6125 0.0000 37.6875 0.5100 ;
    END
  END uart_master.prdata[3]
  PIN uart_master.prdata[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1.1175 39.4800 1.1925 39.9000 ;
    END
  END uart_master.prdata[2]
  PIN uart_master.prdata[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 1.1625 39.3900 1.2375 39.9000 ;
    END
  END uart_master.prdata[1]
  PIN uart_master.prdata[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 37.1625 0.0000 37.2375 0.5100 ;
    END
  END uart_master.prdata[0]
  PIN uart_master.pready
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 37.8675 0.0000 37.9425 0.4200 ;
    END
  END uart_master.pready
  PIN uart_master.pslverr
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 28.8375 0.0000 28.9125 0.4200 ;
    END
  END uart_master.pslverr
  PIN gpio_master.paddr[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 5.6625 40.3200 5.7375 ;
    END
  END gpio_master.paddr[31]
  PIN gpio_master.paddr[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 5.9625 40.3200 6.0375 ;
    END
  END gpio_master.paddr[30]
  PIN gpio_master.paddr[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 6.2625 40.3200 6.3375 ;
    END
  END gpio_master.paddr[29]
  PIN gpio_master.paddr[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 20.3625 39.3900 20.4375 39.9000 ;
    END
  END gpio_master.paddr[28]
  PIN gpio_master.paddr[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 20.6625 39.3900 20.7375 39.9000 ;
    END
  END gpio_master.paddr[27]
  PIN gpio_master.paddr[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 6.5625 40.3200 6.6375 ;
    END
  END gpio_master.paddr[26]
  PIN gpio_master.paddr[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 20.9625 39.3900 21.0375 39.9000 ;
    END
  END gpio_master.paddr[25]
  PIN gpio_master.paddr[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 6.8625 40.3200 6.9375 ;
    END
  END gpio_master.paddr[24]
  PIN gpio_master.paddr[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 7.1625 40.3200 7.2375 ;
    END
  END gpio_master.paddr[23]
  PIN gpio_master.paddr[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 7.4625 40.3200 7.5375 ;
    END
  END gpio_master.paddr[22]
  PIN gpio_master.paddr[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 7.7625 40.3200 7.8375 ;
    END
  END gpio_master.paddr[21]
  PIN gpio_master.paddr[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 21.2625 39.3900 21.3375 39.9000 ;
    END
  END gpio_master.paddr[20]
  PIN gpio_master.paddr[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 8.0625 40.3200 8.1375 ;
    END
  END gpio_master.paddr[19]
  PIN gpio_master.paddr[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 8.3625 40.3200 8.4375 ;
    END
  END gpio_master.paddr[18]
  PIN gpio_master.paddr[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 8.6625 40.3200 8.7375 ;
    END
  END gpio_master.paddr[17]
  PIN gpio_master.paddr[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 8.9625 40.3200 9.0375 ;
    END
  END gpio_master.paddr[16]
  PIN gpio_master.paddr[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 9.2625 40.3200 9.3375 ;
    END
  END gpio_master.paddr[15]
  PIN gpio_master.paddr[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 9.5625 40.3200 9.6375 ;
    END
  END gpio_master.paddr[14]
  PIN gpio_master.paddr[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 9.8625 40.3200 9.9375 ;
    END
  END gpio_master.paddr[13]
  PIN gpio_master.paddr[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 21.5625 39.3900 21.6375 39.9000 ;
    END
  END gpio_master.paddr[12]
  PIN gpio_master.paddr[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 8.2125 39.3900 8.2875 39.9000 ;
    END
  END gpio_master.paddr[11]
  PIN gpio_master.paddr[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 24.7125 0.5100 24.7875 ;
    END
  END gpio_master.paddr[10]
  PIN gpio_master.paddr[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 30.4125 0.5100 30.4875 ;
    END
  END gpio_master.paddr[9]
  PIN gpio_master.paddr[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 14.5125 39.3900 14.5875 39.9000 ;
    END
  END gpio_master.paddr[8]
  PIN gpio_master.paddr[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 27.7125 0.5100 27.7875 ;
    END
  END gpio_master.paddr[7]
  PIN gpio_master.paddr[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 14.2125 39.3900 14.2875 39.9000 ;
    END
  END gpio_master.paddr[6]
  PIN gpio_master.paddr[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 24.7125 0.5100 24.7875 ;
    END
  END gpio_master.paddr[5]
  PIN gpio_master.paddr[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 13.3125 0.5100 13.3875 ;
    END
  END gpio_master.paddr[4]
  PIN gpio_master.paddr[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 28.6125 0.5100 28.6875 ;
    END
  END gpio_master.paddr[3]
  PIN gpio_master.paddr[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 13.9125 39.3900 13.9875 39.9000 ;
    END
  END gpio_master.paddr[2]
  PIN gpio_master.paddr[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12.8775 39.4800 12.9525 39.9000 ;
    END
  END gpio_master.paddr[1]
  PIN gpio_master.paddr[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 9.8625 39.3900 9.9375 39.9000 ;
    END
  END gpio_master.paddr[0]
  PIN gpio_master.pwdata[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 19.0125 0.5100 19.0875 ;
    END
  END gpio_master.pwdata[31]
  PIN gpio_master.pwdata[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 13.3125 0.5100 13.3875 ;
    END
  END gpio_master.pwdata[30]
  PIN gpio_master.pwdata[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 33.1125 0.5100 33.1875 ;
    END
  END gpio_master.pwdata[29]
  PIN gpio_master.pwdata[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 14.5125 0.5100 14.5875 ;
    END
  END gpio_master.pwdata[28]
  PIN gpio_master.pwdata[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18.7125 39.3900 18.7875 39.9000 ;
    END
  END gpio_master.pwdata[27]
  PIN gpio_master.pwdata[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 28.9125 0.5100 28.9875 ;
    END
  END gpio_master.pwdata[26]
  PIN gpio_master.pwdata[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12.7125 39.3900 12.7875 39.9000 ;
    END
  END gpio_master.pwdata[25]
  PIN gpio_master.pwdata[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 20.6475 39.4800 20.7225 39.9000 ;
    END
  END gpio_master.pwdata[24]
  PIN gpio_master.pwdata[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 25.0125 0.5100 25.0875 ;
    END
  END gpio_master.pwdata[23]
  PIN gpio_master.pwdata[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 28.3125 0.5100 28.3875 ;
    END
  END gpio_master.pwdata[22]
  PIN gpio_master.pwdata[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 25.3125 0.5100 25.3875 ;
    END
  END gpio_master.pwdata[21]
  PIN gpio_master.pwdata[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 18.7125 0.5100 18.7875 ;
    END
  END gpio_master.pwdata[20]
  PIN gpio_master.pwdata[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 19.9125 39.3900 19.9875 39.9000 ;
    END
  END gpio_master.pwdata[19]
  PIN gpio_master.pwdata[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4.4625 39.3900 4.5375 39.9000 ;
    END
  END gpio_master.pwdata[18]
  PIN gpio_master.pwdata[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 15.1125 0.5100 15.1875 ;
    END
  END gpio_master.pwdata[17]
  PIN gpio_master.pwdata[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 6.5625 39.3900 6.6375 39.9000 ;
    END
  END gpio_master.pwdata[16]
  PIN gpio_master.pwdata[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 15.5625 39.3900 15.6375 39.9000 ;
    END
  END gpio_master.pwdata[15]
  PIN gpio_master.pwdata[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 15.1125 0.5100 15.1875 ;
    END
  END gpio_master.pwdata[14]
  PIN gpio_master.pwdata[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 14.8125 0.5100 14.8875 ;
    END
  END gpio_master.pwdata[13]
  PIN gpio_master.pwdata[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 26.8125 0.5100 26.8875 ;
    END
  END gpio_master.pwdata[12]
  PIN gpio_master.pwdata[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 13.6125 39.3900 13.6875 39.9000 ;
    END
  END gpio_master.pwdata[11]
  PIN gpio_master.pwdata[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 14.5125 0.5100 14.5875 ;
    END
  END gpio_master.pwdata[10]
  PIN gpio_master.pwdata[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 28.9125 0.5100 28.9875 ;
    END
  END gpio_master.pwdata[9]
  PIN gpio_master.pwdata[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 18.5625 39.3900 18.6375 39.9000 ;
    END
  END gpio_master.pwdata[8]
  PIN gpio_master.pwdata[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 14.8125 0.5100 14.8875 ;
    END
  END gpio_master.pwdata[7]
  PIN gpio_master.pwdata[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12.6675 0.0000 12.7425 0.4200 ;
    END
  END gpio_master.pwdata[6]
  PIN gpio_master.pwdata[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 20.6625 39.3900 20.7375 39.9000 ;
    END
  END gpio_master.pwdata[5]
  PIN gpio_master.pwdata[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 10.9125 0.5100 10.9875 ;
    END
  END gpio_master.pwdata[4]
  PIN gpio_master.pwdata[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 10.9125 0.5100 10.9875 ;
    END
  END gpio_master.pwdata[3]
  PIN gpio_master.pwdata[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 10.6125 0.5100 10.6875 ;
    END
  END gpio_master.pwdata[2]
  PIN gpio_master.pwdata[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 10.6125 0.5100 10.6875 ;
    END
  END gpio_master.pwdata[1]
  PIN gpio_master.pwdata[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11.6625 39.3900 11.7375 39.9000 ;
    END
  END gpio_master.pwdata[0]
  PIN gpio_master.pwrite
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3.8475 0.0000 3.9225 0.4200 ;
    END
  END gpio_master.pwrite
  PIN gpio_master.psel
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 21.4875 39.4800 21.5625 39.9000 ;
    END
  END gpio_master.psel
  PIN gpio_master.penable
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 3.7125 0.5100 3.7875 ;
    END
  END gpio_master.penable
  PIN gpio_master.prdata[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 21.8625 39.3900 21.9375 39.9000 ;
    END
  END gpio_master.prdata[31]
  PIN gpio_master.prdata[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 24.1125 39.3900 24.1875 39.9000 ;
    END
  END gpio_master.prdata[30]
  PIN gpio_master.prdata[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.8100 32.3625 40.3200 32.4375 ;
    END
  END gpio_master.prdata[29]
  PIN gpio_master.prdata[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.8100 10.0125 40.3200 10.0875 ;
    END
  END gpio_master.prdata[28]
  PIN gpio_master.prdata[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.8100 9.7125 40.3200 9.7875 ;
    END
  END gpio_master.prdata[27]
  PIN gpio_master.prdata[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 22.6125 39.3900 22.6875 39.9000 ;
    END
  END gpio_master.prdata[26]
  PIN gpio_master.prdata[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 27.7125 39.3900 27.7875 39.9000 ;
    END
  END gpio_master.prdata[25]
  PIN gpio_master.prdata[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 26.8125 39.3900 26.8875 39.9000 ;
    END
  END gpio_master.prdata[24]
  PIN gpio_master.prdata[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 29.0625 39.3900 29.1375 39.9000 ;
    END
  END gpio_master.prdata[23]
  PIN gpio_master.prdata[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.8100 32.6625 40.3200 32.7375 ;
    END
  END gpio_master.prdata[22]
  PIN gpio_master.prdata[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.8100 9.4125 40.3200 9.4875 ;
    END
  END gpio_master.prdata[21]
  PIN gpio_master.prdata[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.8100 32.9625 40.3200 33.0375 ;
    END
  END gpio_master.prdata[20]
  PIN gpio_master.prdata[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.8100 33.5625 40.3200 33.6375 ;
    END
  END gpio_master.prdata[19]
  PIN gpio_master.prdata[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 38.1975 33.3000 40.3200 33.9000 ;
    END
  END gpio_master.prdata[18]
  PIN gpio_master.prdata[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 25.3125 39.3900 25.3875 39.9000 ;
    END
  END gpio_master.prdata[17]
  PIN gpio_master.prdata[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 25.0125 39.3900 25.0875 39.9000 ;
    END
  END gpio_master.prdata[16]
  PIN gpio_master.prdata[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 23.8125 39.3900 23.8875 39.9000 ;
    END
  END gpio_master.prdata[15]
  PIN gpio_master.prdata[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 20.4375 0.0000 20.5125 0.4200 ;
    END
  END gpio_master.prdata[14]
  PIN gpio_master.prdata[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.8100 9.1125 40.3200 9.1875 ;
    END
  END gpio_master.prdata[13]
  PIN gpio_master.prdata[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 31.9125 39.3900 31.9875 39.9000 ;
    END
  END gpio_master.prdata[12]
  PIN gpio_master.prdata[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 28.6125 39.3900 28.6875 39.9000 ;
    END
  END gpio_master.prdata[11]
  PIN gpio_master.prdata[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 19.4625 39.3900 19.5375 39.9000 ;
    END
  END gpio_master.prdata[10]
  PIN gpio_master.prdata[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.8100 33.8625 40.3200 33.9375 ;
    END
  END gpio_master.prdata[9]
  PIN gpio_master.prdata[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 17.3625 39.3900 17.4375 39.9000 ;
    END
  END gpio_master.prdata[8]
  PIN gpio_master.prdata[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.8100 37.3125 40.3200 37.3875 ;
    END
  END gpio_master.prdata[7]
  PIN gpio_master.prdata[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.8100 34.1625 40.3200 34.2375 ;
    END
  END gpio_master.prdata[6]
  PIN gpio_master.prdata[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 23.5125 39.3900 23.5875 39.9000 ;
    END
  END gpio_master.prdata[5]
  PIN gpio_master.prdata[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 26.0625 39.3900 26.1375 39.9000 ;
    END
  END gpio_master.prdata[4]
  PIN gpio_master.prdata[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.8100 34.4625 40.3200 34.5375 ;
    END
  END gpio_master.prdata[3]
  PIN gpio_master.prdata[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 33.4125 39.3900 33.4875 39.9000 ;
    END
  END gpio_master.prdata[2]
  PIN gpio_master.prdata[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 30.3075 39.4800 30.3825 39.9000 ;
    END
  END gpio_master.prdata[1]
  PIN gpio_master.prdata[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.8100 8.8125 40.3200 8.8875 ;
    END
  END gpio_master.prdata[0]
  PIN gpio_master.pready
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.8100 1.9125 40.3200 1.9875 ;
    END
  END gpio_master.pready
  PIN gpio_master.pslverr
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 30.3075 0.0000 30.3825 0.4200 ;
    END
  END gpio_master.pslverr
  PIN spi_master.paddr[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 10.1625 40.3200 10.2375 ;
    END
  END spi_master.paddr[31]
  PIN spi_master.paddr[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 10.4625 40.3200 10.5375 ;
    END
  END spi_master.paddr[30]
  PIN spi_master.paddr[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 10.7625 40.3200 10.8375 ;
    END
  END spi_master.paddr[29]
  PIN spi_master.paddr[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14.0625 0.0000 14.1375 0.5100 ;
    END
  END spi_master.paddr[28]
  PIN spi_master.paddr[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14.3625 0.0000 14.4375 0.5100 ;
    END
  END spi_master.paddr[27]
  PIN spi_master.paddr[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 11.0625 40.3200 11.1375 ;
    END
  END spi_master.paddr[26]
  PIN spi_master.paddr[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14.6625 0.0000 14.7375 0.5100 ;
    END
  END spi_master.paddr[25]
  PIN spi_master.paddr[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 11.3625 40.3200 11.4375 ;
    END
  END spi_master.paddr[24]
  PIN spi_master.paddr[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 11.6625 40.3200 11.7375 ;
    END
  END spi_master.paddr[23]
  PIN spi_master.paddr[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 11.9625 40.3200 12.0375 ;
    END
  END spi_master.paddr[22]
  PIN spi_master.paddr[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 12.2625 40.3200 12.3375 ;
    END
  END spi_master.paddr[21]
  PIN spi_master.paddr[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14.9625 0.0000 15.0375 0.5100 ;
    END
  END spi_master.paddr[20]
  PIN spi_master.paddr[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 12.5625 40.3200 12.6375 ;
    END
  END spi_master.paddr[19]
  PIN spi_master.paddr[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 12.8625 40.3200 12.9375 ;
    END
  END spi_master.paddr[18]
  PIN spi_master.paddr[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 13.1625 40.3200 13.2375 ;
    END
  END spi_master.paddr[17]
  PIN spi_master.paddr[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 13.4625 40.3200 13.5375 ;
    END
  END spi_master.paddr[16]
  PIN spi_master.paddr[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 13.7625 40.3200 13.8375 ;
    END
  END spi_master.paddr[15]
  PIN spi_master.paddr[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 14.0625 40.3200 14.1375 ;
    END
  END spi_master.paddr[14]
  PIN spi_master.paddr[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15.2625 0.0000 15.3375 0.5100 ;
    END
  END spi_master.paddr[13]
  PIN spi_master.paddr[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 14.3625 40.3200 14.4375 ;
    END
  END spi_master.paddr[12]
  PIN spi_master.paddr[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6.8625 39.3900 6.9375 39.9000 ;
    END
  END spi_master.paddr[11]
  PIN spi_master.paddr[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 6.2625 39.3900 6.3375 39.9000 ;
    END
  END spi_master.paddr[10]
  PIN spi_master.paddr[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 33.7125 0.5100 33.7875 ;
    END
  END spi_master.paddr[9]
  PIN spi_master.paddr[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 5.9625 39.3900 6.0375 39.9000 ;
    END
  END spi_master.paddr[8]
  PIN spi_master.paddr[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 34.0125 0.5100 34.0875 ;
    END
  END spi_master.paddr[7]
  PIN spi_master.paddr[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5.8125 39.3900 5.8875 39.9000 ;
    END
  END spi_master.paddr[6]
  PIN spi_master.paddr[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 5.6625 39.3900 5.7375 39.9000 ;
    END
  END spi_master.paddr[5]
  PIN spi_master.paddr[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 7.9125 0.5100 7.9875 ;
    END
  END spi_master.paddr[4]
  PIN spi_master.paddr[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 34.6125 0.5100 34.6875 ;
    END
  END spi_master.paddr[3]
  PIN spi_master.paddr[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5.5125 39.3900 5.5875 39.9000 ;
    END
  END spi_master.paddr[2]
  PIN spi_master.paddr[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 5.3625 39.3900 5.4375 39.9000 ;
    END
  END spi_master.paddr[1]
  PIN spi_master.paddr[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5.2125 39.3900 5.2875 39.9000 ;
    END
  END spi_master.paddr[0]
  PIN spi_master.pwdata[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 16.0125 0.0000 16.0875 0.5100 ;
    END
  END spi_master.pwdata[31]
  PIN spi_master.pwdata[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11.3625 0.0000 11.4375 0.5100 ;
    END
  END spi_master.pwdata[30]
  PIN spi_master.pwdata[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 34.9125 0.5100 34.9875 ;
    END
  END spi_master.pwdata[29]
  PIN spi_master.pwdata[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 7.6125 0.5100 7.6875 ;
    END
  END spi_master.pwdata[28]
  PIN spi_master.pwdata[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4.9125 39.3900 4.9875 39.9000 ;
    END
  END spi_master.pwdata[27]
  PIN spi_master.pwdata[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 4.7625 39.3900 4.8375 39.9000 ;
    END
  END spi_master.pwdata[26]
  PIN spi_master.pwdata[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 35.2125 0.5100 35.2875 ;
    END
  END spi_master.pwdata[25]
  PIN spi_master.pwdata[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 34.6125 39.3900 34.6875 39.9000 ;
    END
  END spi_master.pwdata[24]
  PIN spi_master.pwdata[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 35.2125 0.5100 35.2875 ;
    END
  END spi_master.pwdata[23]
  PIN spi_master.pwdata[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 4.4625 39.3900 4.5375 39.9000 ;
    END
  END spi_master.pwdata[22]
  PIN spi_master.pwdata[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 35.5125 0.5100 35.5875 ;
    END
  END spi_master.pwdata[21]
  PIN spi_master.pwdata[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 35.5125 0.5100 35.5875 ;
    END
  END spi_master.pwdata[20]
  PIN spi_master.pwdata[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17.7075 0.0000 17.7825 0.4200 ;
    END
  END spi_master.pwdata[19]
  PIN spi_master.pwdata[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3.6375 39.4800 3.7125 39.9000 ;
    END
  END spi_master.pwdata[18]
  PIN spi_master.pwdata[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 7.6125 0.5100 7.6875 ;
    END
  END spi_master.pwdata[17]
  PIN spi_master.pwdata[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 4.1625 39.3900 4.2375 39.9000 ;
    END
  END spi_master.pwdata[16]
  PIN spi_master.pwdata[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 16.7625 0.0000 16.8375 0.5100 ;
    END
  END spi_master.pwdata[15]
  PIN spi_master.pwdata[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 10.9125 0.0000 10.9875 0.5100 ;
    END
  END spi_master.pwdata[14]
  PIN spi_master.pwdata[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 15.4125 0.0000 15.4875 0.5100 ;
    END
  END spi_master.pwdata[13]
  PIN spi_master.pwdata[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 35.8125 0.5100 35.8875 ;
    END
  END spi_master.pwdata[12]
  PIN spi_master.pwdata[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13.2975 0.0000 13.3725 0.4200 ;
    END
  END spi_master.pwdata[11]
  PIN spi_master.pwdata[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 7.3125 0.5100 7.3875 ;
    END
  END spi_master.pwdata[10]
  PIN spi_master.pwdata[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 35.8125 0.5100 35.8875 ;
    END
  END spi_master.pwdata[9]
  PIN spi_master.pwdata[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 3.8625 39.3900 3.9375 39.9000 ;
    END
  END spi_master.pwdata[8]
  PIN spi_master.pwdata[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 7.3125 0.5100 7.3875 ;
    END
  END spi_master.pwdata[7]
  PIN spi_master.pwdata[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15.5625 0.0000 15.6375 0.5100 ;
    END
  END spi_master.pwdata[6]
  PIN spi_master.pwdata[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 18.1125 0.0000 18.1875 0.5100 ;
    END
  END spi_master.pwdata[5]
  PIN spi_master.pwdata[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 10.1625 0.0000 10.2375 0.5100 ;
    END
  END spi_master.pwdata[4]
  PIN spi_master.pwdata[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 0.0000 6.9000 2.1225 7.5000 ;
    END
  END spi_master.pwdata[3]
  PIN spi_master.pwdata[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 7.0125 0.5100 7.0875 ;
    END
  END spi_master.pwdata[2]
  PIN spi_master.pwdata[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 7.0125 0.5100 7.0875 ;
    END
  END spi_master.pwdata[1]
  PIN spi_master.pwdata[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 36.1125 0.5100 36.1875 ;
    END
  END spi_master.pwdata[0]
  PIN spi_master.pwrite
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 3.7125 0.5100 3.7875 ;
    END
  END spi_master.pwrite
  PIN spi_master.psel
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15.1875 0.0000 15.2625 0.4200 ;
    END
  END spi_master.psel
  PIN spi_master.penable
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 3.4125 0.5100 3.4875 ;
    END
  END spi_master.penable
  PIN spi_master.prdata[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 32.8125 39.3900 32.8875 39.9000 ;
    END
  END spi_master.prdata[31]
  PIN spi_master.prdata[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 32.9625 39.3900 33.0375 39.9000 ;
    END
  END spi_master.prdata[30]
  PIN spi_master.prdata[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.8100 37.9125 40.3200 37.9875 ;
    END
  END spi_master.prdata[29]
  PIN spi_master.prdata[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.8100 4.6125 40.3200 4.6875 ;
    END
  END spi_master.prdata[28]
  PIN spi_master.prdata[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.8100 4.3125 40.3200 4.3875 ;
    END
  END spi_master.prdata[27]
  PIN spi_master.prdata[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 33.1125 39.3900 33.1875 39.9000 ;
    END
  END spi_master.prdata[26]
  PIN spi_master.prdata[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 33.4125 39.3900 33.4875 39.9000 ;
    END
  END spi_master.prdata[25]
  PIN spi_master.prdata[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 33.7125 39.3900 33.7875 39.9000 ;
    END
  END spi_master.prdata[24]
  PIN spi_master.prdata[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 34.0125 39.3900 34.0875 39.9000 ;
    END
  END spi_master.prdata[23]
  PIN spi_master.prdata[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.8100 38.2125 40.3200 38.2875 ;
    END
  END spi_master.prdata[22]
  PIN spi_master.prdata[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.8100 4.0125 40.3200 4.0875 ;
    END
  END spi_master.prdata[21]
  PIN spi_master.prdata[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.8100 38.5125 40.3200 38.5875 ;
    END
  END spi_master.prdata[20]
  PIN spi_master.prdata[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 38.9175 39.4800 38.9925 39.9000 ;
    END
  END spi_master.prdata[19]
  PIN spi_master.prdata[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.8100 38.8125 40.3200 38.8875 ;
    END
  END spi_master.prdata[18]
  PIN spi_master.prdata[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 25.4625 0.0000 25.5375 0.5100 ;
    END
  END spi_master.prdata[17]
  PIN spi_master.prdata[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 24.2625 0.0000 24.3375 0.5100 ;
    END
  END spi_master.prdata[16]
  PIN spi_master.prdata[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 23.9625 0.0000 24.0375 0.5100 ;
    END
  END spi_master.prdata[15]
  PIN spi_master.prdata[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 19.4625 0.0000 19.5375 0.5100 ;
    END
  END spi_master.prdata[14]
  PIN spi_master.prdata[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.8100 3.7125 40.3200 3.7875 ;
    END
  END spi_master.prdata[13]
  PIN spi_master.prdata[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 34.0125 39.3900 34.0875 39.9000 ;
    END
  END spi_master.prdata[12]
  PIN spi_master.prdata[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 29.2125 0.0000 29.2875 0.5100 ;
    END
  END spi_master.prdata[11]
  PIN spi_master.prdata[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 34.6125 0.5100 34.6875 ;
    END
  END spi_master.prdata[10]
  PIN spi_master.prdata[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 39.2625 39.3900 39.3375 39.9000 ;
    END
  END spi_master.prdata[9]
  PIN spi_master.prdata[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 5.0625 39.3900 5.1375 39.9000 ;
    END
  END spi_master.prdata[8]
  PIN spi_master.prdata[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 38.4975 39.4800 38.5725 39.9000 ;
    END
  END spi_master.prdata[7]
  PIN spi_master.prdata[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 39.4125 39.3900 39.4875 39.9000 ;
    END
  END spi_master.prdata[6]
  PIN spi_master.prdata[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 22.9575 0.0000 23.0325 0.4200 ;
    END
  END spi_master.prdata[5]
  PIN spi_master.prdata[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 34.3125 39.3900 34.3875 39.9000 ;
    END
  END spi_master.prdata[4]
  PIN spi_master.prdata[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 38.9625 39.3900 39.0375 39.9000 ;
    END
  END spi_master.prdata[3]
  PIN spi_master.prdata[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 34.3125 39.3900 34.3875 39.9000 ;
    END
  END spi_master.prdata[2]
  PIN spi_master.prdata[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 34.7175 39.4800 34.7925 39.9000 ;
    END
  END spi_master.prdata[1]
  PIN spi_master.prdata[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.8100 3.4125 40.3200 3.4875 ;
    END
  END spi_master.prdata[0]
  PIN spi_master.pready
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.8100 1.6125 40.3200 1.6875 ;
    END
  END spi_master.pready
  PIN spi_master.pslverr
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 31.1625 0.0000 31.2375 0.5100 ;
    END
  END spi_master.pslverr
  PIN timer_master.paddr[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 14.6625 40.3200 14.7375 ;
    END
  END timer_master.paddr[31]
  PIN timer_master.paddr[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 14.9625 40.3200 15.0375 ;
    END
  END timer_master.paddr[30]
  PIN timer_master.paddr[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 15.2625 40.3200 15.3375 ;
    END
  END timer_master.paddr[29]
  PIN timer_master.paddr[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 18.4125 0.0000 18.4875 0.5100 ;
    END
  END timer_master.paddr[28]
  PIN timer_master.paddr[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 18.7125 0.0000 18.7875 0.5100 ;
    END
  END timer_master.paddr[27]
  PIN timer_master.paddr[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 15.5625 40.3200 15.6375 ;
    END
  END timer_master.paddr[26]
  PIN timer_master.paddr[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18.7125 0.0000 18.7875 0.5100 ;
    END
  END timer_master.paddr[25]
  PIN timer_master.paddr[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 15.8625 40.3200 15.9375 ;
    END
  END timer_master.paddr[24]
  PIN timer_master.paddr[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 16.1625 40.3200 16.2375 ;
    END
  END timer_master.paddr[23]
  PIN timer_master.paddr[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 16.4625 40.3200 16.5375 ;
    END
  END timer_master.paddr[22]
  PIN timer_master.paddr[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 16.7625 40.3200 16.8375 ;
    END
  END timer_master.paddr[21]
  PIN timer_master.paddr[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 19.0125 0.0000 19.0875 0.5100 ;
    END
  END timer_master.paddr[20]
  PIN timer_master.paddr[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 17.0625 40.3200 17.1375 ;
    END
  END timer_master.paddr[19]
  PIN timer_master.paddr[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 17.3625 40.3200 17.4375 ;
    END
  END timer_master.paddr[18]
  PIN timer_master.paddr[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 17.6625 40.3200 17.7375 ;
    END
  END timer_master.paddr[17]
  PIN timer_master.paddr[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 17.9625 40.3200 18.0375 ;
    END
  END timer_master.paddr[16]
  PIN timer_master.paddr[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 18.2625 40.3200 18.3375 ;
    END
  END timer_master.paddr[15]
  PIN timer_master.paddr[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 18.5625 40.3200 18.6375 ;
    END
  END timer_master.paddr[14]
  PIN timer_master.paddr[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 19.3125 0.0000 19.3875 0.5100 ;
    END
  END timer_master.paddr[13]
  PIN timer_master.paddr[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 19.6125 0.0000 19.6875 0.5100 ;
    END
  END timer_master.paddr[12]
  PIN timer_master.paddr[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3.7125 39.3900 3.7875 39.9000 ;
    END
  END timer_master.paddr[11]
  PIN timer_master.paddr[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9.1125 0.0000 9.1875 0.5100 ;
    END
  END timer_master.paddr[10]
  PIN timer_master.paddr[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 36.1125 0.5100 36.1875 ;
    END
  END timer_master.paddr[9]
  PIN timer_master.paddr[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 3.5625 39.3900 3.6375 39.9000 ;
    END
  END timer_master.paddr[8]
  PIN timer_master.paddr[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 36.4125 0.5100 36.4875 ;
    END
  END timer_master.paddr[7]
  PIN timer_master.paddr[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3.4125 39.3900 3.4875 39.9000 ;
    END
  END timer_master.paddr[6]
  PIN timer_master.paddr[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 11.3625 0.0000 11.4375 0.5100 ;
    END
  END timer_master.paddr[5]
  PIN timer_master.paddr[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8.4675 0.0000 8.5425 0.4200 ;
    END
  END timer_master.paddr[4]
  PIN timer_master.paddr[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3.2175 39.4800 3.2925 39.9000 ;
    END
  END timer_master.paddr[3]
  PIN timer_master.paddr[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 3.2625 39.3900 3.3375 39.9000 ;
    END
  END timer_master.paddr[2]
  PIN timer_master.paddr[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 36.7125 0.5100 36.7875 ;
    END
  END timer_master.paddr[1]
  PIN timer_master.paddr[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 36.7125 0.5100 36.7875 ;
    END
  END timer_master.paddr[0]
  PIN timer_master.pwdata[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 14.9625 0.0000 15.0375 0.5100 ;
    END
  END timer_master.pwdata[31]
  PIN timer_master.pwdata[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10.5675 0.0000 10.6425 0.4200 ;
    END
  END timer_master.pwdata[30]
  PIN timer_master.pwdata[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 2.9625 39.3900 3.0375 39.9000 ;
    END
  END timer_master.pwdata[29]
  PIN timer_master.pwdata[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 6.7125 0.5100 6.7875 ;
    END
  END timer_master.pwdata[28]
  PIN timer_master.pwdata[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 37.0125 0.5100 37.0875 ;
    END
  END timer_master.pwdata[27]
  PIN timer_master.pwdata[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 37.0125 0.5100 37.0875 ;
    END
  END timer_master.pwdata[26]
  PIN timer_master.pwdata[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2.8125 39.3900 2.8875 39.9000 ;
    END
  END timer_master.pwdata[25]
  PIN timer_master.pwdata[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 2.6625 39.3900 2.7375 39.9000 ;
    END
  END timer_master.pwdata[24]
  PIN timer_master.pwdata[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 37.3125 0.5100 37.3875 ;
    END
  END timer_master.pwdata[23]
  PIN timer_master.pwdata[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 37.3125 0.5100 37.3875 ;
    END
  END timer_master.pwdata[22]
  PIN timer_master.pwdata[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2.5125 39.3900 2.5875 39.9000 ;
    END
  END timer_master.pwdata[21]
  PIN timer_master.pwdata[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2.3775 39.4800 2.4525 39.9000 ;
    END
  END timer_master.pwdata[20]
  PIN timer_master.pwdata[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 17.6625 0.0000 17.7375 0.5100 ;
    END
  END timer_master.pwdata[19]
  PIN timer_master.pwdata[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 2.3625 39.3900 2.4375 39.9000 ;
    END
  END timer_master.pwdata[18]
  PIN timer_master.pwdata[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 6.7125 0.5100 6.7875 ;
    END
  END timer_master.pwdata[17]
  PIN timer_master.pwdata[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 37.6125 0.5100 37.6875 ;
    END
  END timer_master.pwdata[16]
  PIN timer_master.pwdata[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16.6125 0.0000 16.6875 0.5100 ;
    END
  END timer_master.pwdata[15]
  PIN timer_master.pwdata[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10.6125 0.0000 10.6875 0.5100 ;
    END
  END timer_master.pwdata[14]
  PIN timer_master.pwdata[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 13.3125 0.0000 13.3875 0.5100 ;
    END
  END timer_master.pwdata[13]
  PIN timer_master.pwdata[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 6.4125 0.5100 6.4875 ;
    END
  END timer_master.pwdata[12]
  PIN timer_master.pwdata[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14.7675 0.0000 14.8425 0.4200 ;
    END
  END timer_master.pwdata[11]
  PIN timer_master.pwdata[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 6.4125 0.5100 6.4875 ;
    END
  END timer_master.pwdata[10]
  PIN timer_master.pwdata[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 37.6125 0.5100 37.6875 ;
    END
  END timer_master.pwdata[9]
  PIN timer_master.pwdata[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2.2125 39.3900 2.2875 39.9000 ;
    END
  END timer_master.pwdata[8]
  PIN timer_master.pwdata[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6.1575 0.0000 6.2325 0.4200 ;
    END
  END timer_master.pwdata[7]
  PIN timer_master.pwdata[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 14.6625 0.0000 14.7375 0.5100 ;
    END
  END timer_master.pwdata[6]
  PIN timer_master.pwdata[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 20.0625 0.0000 20.1375 0.5100 ;
    END
  END timer_master.pwdata[5]
  PIN timer_master.pwdata[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9.8625 0.0000 9.9375 0.5100 ;
    END
  END timer_master.pwdata[4]
  PIN timer_master.pwdata[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 6.1125 0.5100 6.1875 ;
    END
  END timer_master.pwdata[3]
  PIN timer_master.pwdata[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 6.1125 0.5100 6.1875 ;
    END
  END timer_master.pwdata[2]
  PIN timer_master.pwdata[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 5.8125 0.5100 5.8875 ;
    END
  END timer_master.pwdata[1]
  PIN timer_master.pwdata[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 2.0625 39.3900 2.1375 39.9000 ;
    END
  END timer_master.pwdata[0]
  PIN timer_master.pwrite
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3.4275 0.0000 3.5025 0.4200 ;
    END
  END timer_master.pwrite
  PIN timer_master.psel
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 19.5975 0.0000 19.6725 0.4200 ;
    END
  END timer_master.psel
  PIN timer_master.penable
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 3.4125 0.5100 3.4875 ;
    END
  END timer_master.penable
  PIN timer_master.prdata[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 34.6125 39.3900 34.6875 39.9000 ;
    END
  END timer_master.prdata[31]
  PIN timer_master.prdata[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 34.9125 39.3900 34.9875 39.9000 ;
    END
  END timer_master.prdata[30]
  PIN timer_master.prdata[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 37.4625 39.3900 37.5375 39.9000 ;
    END
  END timer_master.prdata[29]
  PIN timer_master.prdata[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 36.3975 0.0000 36.4725 0.4200 ;
    END
  END timer_master.prdata[28]
  PIN timer_master.prdata[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 36.8175 0.0000 36.8925 0.4200 ;
    END
  END timer_master.prdata[27]
  PIN timer_master.prdata[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 34.9125 39.3900 34.9875 39.9000 ;
    END
  END timer_master.prdata[26]
  PIN timer_master.prdata[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 35.1375 39.4800 35.2125 39.9000 ;
    END
  END timer_master.prdata[25]
  PIN timer_master.prdata[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 27.5625 0.0000 27.6375 0.5100 ;
    END
  END timer_master.prdata[24]
  PIN timer_master.prdata[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 35.2125 39.3900 35.2875 39.9000 ;
    END
  END timer_master.prdata[23]
  PIN timer_master.prdata[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 37.0125 39.3900 37.0875 39.9000 ;
    END
  END timer_master.prdata[22]
  PIN timer_master.prdata[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.8100 3.1125 40.3200 3.1875 ;
    END
  END timer_master.prdata[21]
  PIN timer_master.prdata[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 37.4625 39.3900 37.5375 39.9000 ;
    END
  END timer_master.prdata[20]
  PIN timer_master.prdata[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 37.6575 39.4800 37.7325 39.9000 ;
    END
  END timer_master.prdata[19]
  PIN timer_master.prdata[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 37.0125 39.3900 37.0875 39.9000 ;
    END
  END timer_master.prdata[18]
  PIN timer_master.prdata[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 26.9475 0.0000 27.0225 0.4200 ;
    END
  END timer_master.prdata[17]
  PIN timer_master.prdata[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 25.6875 0.0000 25.7625 0.4200 ;
    END
  END timer_master.prdata[16]
  PIN timer_master.prdata[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 23.5875 0.0000 23.6625 0.4200 ;
    END
  END timer_master.prdata[15]
  PIN timer_master.prdata[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 20.0175 0.0000 20.0925 0.4200 ;
    END
  END timer_master.prdata[14]
  PIN timer_master.prdata[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.8100 2.8125 40.3200 2.8875 ;
    END
  END timer_master.prdata[13]
  PIN timer_master.prdata[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 35.2125 39.3900 35.2875 39.9000 ;
    END
  END timer_master.prdata[12]
  PIN timer_master.prdata[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 26.6625 0.0000 26.7375 0.5100 ;
    END
  END timer_master.prdata[11]
  PIN timer_master.prdata[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 35.5125 39.3900 35.5875 39.9000 ;
    END
  END timer_master.prdata[10]
  PIN timer_master.prdata[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 35.8125 39.3900 35.8875 39.9000 ;
    END
  END timer_master.prdata[9]
  PIN timer_master.prdata[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3.1125 39.3900 3.1875 39.9000 ;
    END
  END timer_master.prdata[8]
  PIN timer_master.prdata[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 36.1125 39.3900 36.1875 39.9000 ;
    END
  END timer_master.prdata[7]
  PIN timer_master.prdata[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 37.7625 39.3900 37.8375 39.9000 ;
    END
  END timer_master.prdata[6]
  PIN timer_master.prdata[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 22.4625 0.0000 22.5375 0.5100 ;
    END
  END timer_master.prdata[5]
  PIN timer_master.prdata[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 35.5125 39.3900 35.5875 39.9000 ;
    END
  END timer_master.prdata[4]
  PIN timer_master.prdata[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 36.5625 39.3900 36.6375 39.9000 ;
    END
  END timer_master.prdata[3]
  PIN timer_master.prdata[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 36.7125 39.3900 36.7875 39.9000 ;
    END
  END timer_master.prdata[2]
  PIN timer_master.prdata[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 38.0775 39.4800 38.1525 39.9000 ;
    END
  END timer_master.prdata[1]
  PIN timer_master.prdata[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 35.7675 0.0000 35.8425 0.4200 ;
    END
  END timer_master.prdata[0]
  PIN timer_master.pready
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 34.7175 0.0000 34.7925 0.4200 ;
    END
  END timer_master.pready
  PIN timer_master.pslverr
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 31.7625 0.0000 31.8375 0.5100 ;
    END
  END timer_master.pslverr
  PIN event_unit_master.paddr[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 18.8625 40.3200 18.9375 ;
    END
  END event_unit_master.paddr[31]
  PIN event_unit_master.paddr[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 19.1625 40.3200 19.2375 ;
    END
  END event_unit_master.paddr[30]
  PIN event_unit_master.paddr[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 19.4625 40.3200 19.5375 ;
    END
  END event_unit_master.paddr[29]
  PIN event_unit_master.paddr[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15.7125 39.3900 15.7875 39.9000 ;
    END
  END event_unit_master.paddr[28]
  PIN event_unit_master.paddr[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16.0125 39.3900 16.0875 39.9000 ;
    END
  END event_unit_master.paddr[27]
  PIN event_unit_master.paddr[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 19.7625 40.3200 19.8375 ;
    END
  END event_unit_master.paddr[26]
  PIN event_unit_master.paddr[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16.3125 39.3900 16.3875 39.9000 ;
    END
  END event_unit_master.paddr[25]
  PIN event_unit_master.paddr[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 20.0625 40.3200 20.1375 ;
    END
  END event_unit_master.paddr[24]
  PIN event_unit_master.paddr[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 20.3625 40.3200 20.4375 ;
    END
  END event_unit_master.paddr[23]
  PIN event_unit_master.paddr[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 20.6625 40.3200 20.7375 ;
    END
  END event_unit_master.paddr[22]
  PIN event_unit_master.paddr[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 20.9625 40.3200 21.0375 ;
    END
  END event_unit_master.paddr[21]
  PIN event_unit_master.paddr[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16.6125 39.3900 16.6875 39.9000 ;
    END
  END event_unit_master.paddr[20]
  PIN event_unit_master.paddr[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 21.2625 40.3200 21.3375 ;
    END
  END event_unit_master.paddr[19]
  PIN event_unit_master.paddr[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 21.5625 40.3200 21.6375 ;
    END
  END event_unit_master.paddr[18]
  PIN event_unit_master.paddr[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 21.8625 40.3200 21.9375 ;
    END
  END event_unit_master.paddr[17]
  PIN event_unit_master.paddr[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 22.1625 40.3200 22.2375 ;
    END
  END event_unit_master.paddr[16]
  PIN event_unit_master.paddr[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 22.4625 40.3200 22.5375 ;
    END
  END event_unit_master.paddr[15]
  PIN event_unit_master.paddr[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16.9125 39.3900 16.9875 39.9000 ;
    END
  END event_unit_master.paddr[14]
  PIN event_unit_master.paddr[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 22.7625 40.3200 22.8375 ;
    END
  END event_unit_master.paddr[13]
  PIN event_unit_master.paddr[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 23.0625 40.3200 23.1375 ;
    END
  END event_unit_master.paddr[12]
  PIN event_unit_master.paddr[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7.1625 39.3900 7.2375 39.9000 ;
    END
  END event_unit_master.paddr[11]
  PIN event_unit_master.paddr[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 25.9125 0.5100 25.9875 ;
    END
  END event_unit_master.paddr[10]
  PIN event_unit_master.paddr[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7.7625 39.3900 7.8375 39.9000 ;
    END
  END event_unit_master.paddr[9]
  PIN event_unit_master.paddr[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13.4625 39.3900 13.5375 39.9000 ;
    END
  END event_unit_master.paddr[8]
  PIN event_unit_master.paddr[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 25.6125 0.5100 25.6875 ;
    END
  END event_unit_master.paddr[7]
  PIN event_unit_master.paddr[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 16.4625 39.3900 16.5375 39.9000 ;
    END
  END event_unit_master.paddr[6]
  PIN event_unit_master.paddr[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 24.4125 0.5100 24.4875 ;
    END
  END event_unit_master.paddr[5]
  PIN event_unit_master.paddr[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 16.0125 0.5100 16.0875 ;
    END
  END event_unit_master.paddr[4]
  PIN event_unit_master.paddr[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 0.0000 29.7000 2.1225 30.3000 ;
    END
  END event_unit_master.paddr[3]
  PIN event_unit_master.paddr[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17.2875 39.4800 17.3625 39.9000 ;
    END
  END event_unit_master.paddr[2]
  PIN event_unit_master.paddr[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11.3625 39.3900 11.4375 39.9000 ;
    END
  END event_unit_master.paddr[1]
  PIN event_unit_master.paddr[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 9.5625 39.3900 9.6375 39.9000 ;
    END
  END event_unit_master.paddr[0]
  PIN event_unit_master.pwdata[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 20.5125 0.5100 20.5875 ;
    END
  END event_unit_master.pwdata[31]
  PIN event_unit_master.pwdata[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 16.0125 0.5100 16.0875 ;
    END
  END event_unit_master.pwdata[30]
  PIN event_unit_master.pwdata[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 34.3125 0.5100 34.3875 ;
    END
  END event_unit_master.pwdata[29]
  PIN event_unit_master.pwdata[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 15.4125 0.5100 15.4875 ;
    END
  END event_unit_master.pwdata[28]
  PIN event_unit_master.pwdata[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 17.9625 39.3900 18.0375 39.9000 ;
    END
  END event_unit_master.pwdata[27]
  PIN event_unit_master.pwdata[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 32.5125 0.5100 32.5875 ;
    END
  END event_unit_master.pwdata[26]
  PIN event_unit_master.pwdata[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11.1975 39.4800 11.2725 39.9000 ;
    END
  END event_unit_master.pwdata[25]
  PIN event_unit_master.pwdata[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 19.6125 39.3900 19.6875 39.9000 ;
    END
  END event_unit_master.pwdata[24]
  PIN event_unit_master.pwdata[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 24.1125 0.5100 24.1875 ;
    END
  END event_unit_master.pwdata[23]
  PIN event_unit_master.pwdata[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 26.2125 0.5100 26.2875 ;
    END
  END event_unit_master.pwdata[22]
  PIN event_unit_master.pwdata[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 25.6125 0.5100 25.6875 ;
    END
  END event_unit_master.pwdata[21]
  PIN event_unit_master.pwdata[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 20.6625 0.5100 20.7375 ;
    END
  END event_unit_master.pwdata[20]
  PIN event_unit_master.pwdata[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18.9675 0.0000 19.0425 0.4200 ;
    END
  END event_unit_master.pwdata[19]
  PIN event_unit_master.pwdata[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2.7975 39.4800 2.8725 39.9000 ;
    END
  END event_unit_master.pwdata[18]
  PIN event_unit_master.pwdata[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 17.9625 0.5100 18.0375 ;
    END
  END event_unit_master.pwdata[17]
  PIN event_unit_master.pwdata[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4.6875 39.4800 4.7625 39.9000 ;
    END
  END event_unit_master.pwdata[16]
  PIN event_unit_master.pwdata[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16.0275 39.4800 16.1025 39.9000 ;
    END
  END event_unit_master.pwdata[15]
  PIN event_unit_master.pwdata[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 17.8125 0.5100 17.8875 ;
    END
  END event_unit_master.pwdata[14]
  PIN event_unit_master.pwdata[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 0.0000 17.7000 2.1225 18.3000 ;
    END
  END event_unit_master.pwdata[13]
  PIN event_unit_master.pwdata[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 23.5125 0.5100 23.5875 ;
    END
  END event_unit_master.pwdata[12]
  PIN event_unit_master.pwdata[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 14.8125 39.3900 14.8875 39.9000 ;
    END
  END event_unit_master.pwdata[11]
  PIN event_unit_master.pwdata[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 15.7125 0.5100 15.7875 ;
    END
  END event_unit_master.pwdata[10]
  PIN event_unit_master.pwdata[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 26.5125 0.5100 26.5875 ;
    END
  END event_unit_master.pwdata[9]
  PIN event_unit_master.pwdata[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 15.8625 39.3900 15.9375 39.9000 ;
    END
  END event_unit_master.pwdata[8]
  PIN event_unit_master.pwdata[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 16.9125 0.5100 16.9875 ;
    END
  END event_unit_master.pwdata[7]
  PIN event_unit_master.pwdata[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 17.0625 0.0000 17.1375 0.5100 ;
    END
  END event_unit_master.pwdata[6]
  PIN event_unit_master.pwdata[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 18.2625 39.3900 18.3375 39.9000 ;
    END
  END event_unit_master.pwdata[5]
  PIN event_unit_master.pwdata[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 16.3125 0.5100 16.3875 ;
    END
  END event_unit_master.pwdata[4]
  PIN event_unit_master.pwdata[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 15.7125 0.5100 15.7875 ;
    END
  END event_unit_master.pwdata[3]
  PIN event_unit_master.pwdata[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 16.7625 0.5100 16.8375 ;
    END
  END event_unit_master.pwdata[2]
  PIN event_unit_master.pwdata[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 16.3125 0.5100 16.3875 ;
    END
  END event_unit_master.pwdata[1]
  PIN event_unit_master.pwdata[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 24.1125 0.5100 24.1875 ;
    END
  END event_unit_master.pwdata[0]
  PIN event_unit_master.pwrite
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 3.1125 0.5100 3.1875 ;
    END
  END event_unit_master.pwrite
  PIN event_unit_master.psel
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16.8675 39.4800 16.9425 39.9000 ;
    END
  END event_unit_master.psel
  PIN event_unit_master.penable
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 2.8125 0.5100 2.8875 ;
    END
  END event_unit_master.penable
  PIN event_unit_master.prdata[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 21.0675 39.4800 21.1425 39.9000 ;
    END
  END event_unit_master.prdata[31]
  PIN event_unit_master.prdata[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 24.4125 39.3900 24.4875 39.9000 ;
    END
  END event_unit_master.prdata[30]
  PIN event_unit_master.prdata[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.8100 29.9625 40.3200 30.0375 ;
    END
  END event_unit_master.prdata[29]
  PIN event_unit_master.prdata[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.8100 19.7625 40.3200 19.8375 ;
    END
  END event_unit_master.prdata[28]
  PIN event_unit_master.prdata[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.8100 15.5625 40.3200 15.6375 ;
    END
  END event_unit_master.prdata[27]
  PIN event_unit_master.prdata[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 23.2125 39.3900 23.2875 39.9000 ;
    END
  END event_unit_master.prdata[26]
  PIN event_unit_master.prdata[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 27.1125 39.3900 27.1875 39.9000 ;
    END
  END event_unit_master.prdata[25]
  PIN event_unit_master.prdata[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.8100 26.6625 40.3200 26.7375 ;
    END
  END event_unit_master.prdata[24]
  PIN event_unit_master.prdata[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.8100 26.3625 40.3200 26.4375 ;
    END
  END event_unit_master.prdata[23]
  PIN event_unit_master.prdata[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.8100 26.9625 40.3200 27.0375 ;
    END
  END event_unit_master.prdata[22]
  PIN event_unit_master.prdata[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.8100 17.6625 40.3200 17.7375 ;
    END
  END event_unit_master.prdata[21]
  PIN event_unit_master.prdata[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 38.1975 28.5000 40.3200 29.1000 ;
    END
  END event_unit_master.prdata[20]
  PIN event_unit_master.prdata[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.8100 32.0625 40.3200 32.1375 ;
    END
  END event_unit_master.prdata[19]
  PIN event_unit_master.prdata[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.8100 22.4625 40.3200 22.5375 ;
    END
  END event_unit_master.prdata[18]
  PIN event_unit_master.prdata[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.8100 18.8625 40.3200 18.9375 ;
    END
  END event_unit_master.prdata[17]
  PIN event_unit_master.prdata[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 25.6125 39.3900 25.6875 39.9000 ;
    END
  END event_unit_master.prdata[16]
  PIN event_unit_master.prdata[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.8100 20.0625 40.3200 20.1375 ;
    END
  END event_unit_master.prdata[15]
  PIN event_unit_master.prdata[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.8100 18.5625 40.3200 18.6375 ;
    END
  END event_unit_master.prdata[14]
  PIN event_unit_master.prdata[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.8100 14.5125 40.3200 14.5875 ;
    END
  END event_unit_master.prdata[13]
  PIN event_unit_master.prdata[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 31.3575 39.4800 31.4325 39.9000 ;
    END
  END event_unit_master.prdata[12]
  PIN event_unit_master.prdata[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.8100 22.1625 40.3200 22.2375 ;
    END
  END event_unit_master.prdata[11]
  PIN event_unit_master.prdata[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 19.1625 39.3900 19.2375 39.9000 ;
    END
  END event_unit_master.prdata[10]
  PIN event_unit_master.prdata[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.8100 21.8625 40.3200 21.9375 ;
    END
  END event_unit_master.prdata[9]
  PIN event_unit_master.prdata[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17.6625 39.3900 17.7375 39.9000 ;
    END
  END event_unit_master.prdata[8]
  PIN event_unit_master.prdata[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 32.8275 39.4800 32.9025 39.9000 ;
    END
  END event_unit_master.prdata[7]
  PIN event_unit_master.prdata[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.8100 23.8125 40.3200 23.8875 ;
    END
  END event_unit_master.prdata[6]
  PIN event_unit_master.prdata[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 22.1175 39.4800 22.1925 39.9000 ;
    END
  END event_unit_master.prdata[5]
  PIN event_unit_master.prdata[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 25.3125 39.3900 25.3875 39.9000 ;
    END
  END event_unit_master.prdata[4]
  PIN event_unit_master.prdata[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 38.1975 24.9000 40.3200 25.5000 ;
    END
  END event_unit_master.prdata[3]
  PIN event_unit_master.prdata[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 28.7625 39.3900 28.8375 39.9000 ;
    END
  END event_unit_master.prdata[2]
  PIN event_unit_master.prdata[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 29.8125 39.3900 29.8875 39.9000 ;
    END
  END event_unit_master.prdata[1]
  PIN event_unit_master.prdata[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 38.1975 15.3000 40.3200 15.9000 ;
    END
  END event_unit_master.prdata[0]
  PIN event_unit_master.pready
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 34.0125 0.0000 34.0875 0.5100 ;
    END
  END event_unit_master.pready
  PIN event_unit_master.pslverr
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 31.7625 0.0000 31.8375 0.5100 ;
    END
  END event_unit_master.pslverr
  PIN i2c_master.paddr[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 23.3625 40.3200 23.4375 ;
    END
  END i2c_master.paddr[31]
  PIN i2c_master.paddr[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 23.6625 40.3200 23.7375 ;
    END
  END i2c_master.paddr[30]
  PIN i2c_master.paddr[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 23.9625 40.3200 24.0375 ;
    END
  END i2c_master.paddr[29]
  PIN i2c_master.paddr[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 20.0625 0.0000 20.1375 0.5100 ;
    END
  END i2c_master.paddr[28]
  PIN i2c_master.paddr[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 20.3625 0.0000 20.4375 0.5100 ;
    END
  END i2c_master.paddr[27]
  PIN i2c_master.paddr[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 24.2625 40.3200 24.3375 ;
    END
  END i2c_master.paddr[26]
  PIN i2c_master.paddr[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 20.6625 0.0000 20.7375 0.5100 ;
    END
  END i2c_master.paddr[25]
  PIN i2c_master.paddr[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 24.5625 40.3200 24.6375 ;
    END
  END i2c_master.paddr[24]
  PIN i2c_master.paddr[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 24.8625 40.3200 24.9375 ;
    END
  END i2c_master.paddr[23]
  PIN i2c_master.paddr[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 25.1625 40.3200 25.2375 ;
    END
  END i2c_master.paddr[22]
  PIN i2c_master.paddr[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 25.4625 40.3200 25.5375 ;
    END
  END i2c_master.paddr[21]
  PIN i2c_master.paddr[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 20.9625 0.0000 21.0375 0.5100 ;
    END
  END i2c_master.paddr[20]
  PIN i2c_master.paddr[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 25.7625 40.3200 25.8375 ;
    END
  END i2c_master.paddr[19]
  PIN i2c_master.paddr[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 26.0625 40.3200 26.1375 ;
    END
  END i2c_master.paddr[18]
  PIN i2c_master.paddr[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 26.3625 40.3200 26.4375 ;
    END
  END i2c_master.paddr[17]
  PIN i2c_master.paddr[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 26.6625 40.3200 26.7375 ;
    END
  END i2c_master.paddr[16]
  PIN i2c_master.paddr[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 26.9625 40.3200 27.0375 ;
    END
  END i2c_master.paddr[15]
  PIN i2c_master.paddr[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 21.2625 0.0000 21.3375 0.5100 ;
    END
  END i2c_master.paddr[14]
  PIN i2c_master.paddr[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 27.2625 40.3200 27.3375 ;
    END
  END i2c_master.paddr[13]
  PIN i2c_master.paddr[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 21.5625 0.0000 21.6375 0.5100 ;
    END
  END i2c_master.paddr[12]
  PIN i2c_master.paddr[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8.4675 39.4800 8.5425 39.9000 ;
    END
  END i2c_master.paddr[11]
  PIN i2c_master.paddr[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 29.2125 0.5100 29.2875 ;
    END
  END i2c_master.paddr[10]
  PIN i2c_master.paddr[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 10.3125 39.3900 10.3875 39.9000 ;
    END
  END i2c_master.paddr[9]
  PIN i2c_master.paddr[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 15.1125 39.3900 15.1875 39.9000 ;
    END
  END i2c_master.paddr[8]
  PIN i2c_master.paddr[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 29.5125 0.5100 29.5875 ;
    END
  END i2c_master.paddr[7]
  PIN i2c_master.paddr[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 13.3125 39.3900 13.3875 39.9000 ;
    END
  END i2c_master.paddr[6]
  PIN i2c_master.paddr[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10.5675 39.4800 10.6425 39.9000 ;
    END
  END i2c_master.paddr[5]
  PIN i2c_master.paddr[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 10.3125 0.5100 10.3875 ;
    END
  END i2c_master.paddr[4]
  PIN i2c_master.paddr[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 29.8125 0.5100 29.8875 ;
    END
  END i2c_master.paddr[3]
  PIN i2c_master.paddr[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13.1625 39.3900 13.2375 39.9000 ;
    END
  END i2c_master.paddr[2]
  PIN i2c_master.paddr[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 11.6625 39.3900 11.7375 39.9000 ;
    END
  END i2c_master.paddr[1]
  PIN i2c_master.paddr[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9.2625 39.3900 9.3375 39.9000 ;
    END
  END i2c_master.paddr[0]
  PIN i2c_master.pwdata[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13.7625 0.0000 13.8375 0.5100 ;
    END
  END i2c_master.pwdata[31]
  PIN i2c_master.pwdata[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12.4125 0.0000 12.4875 0.5100 ;
    END
  END i2c_master.pwdata[30]
  PIN i2c_master.pwdata[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 32.2125 0.5100 32.2875 ;
    END
  END i2c_master.pwdata[29]
  PIN i2c_master.pwdata[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 10.3125 0.5100 10.3875 ;
    END
  END i2c_master.pwdata[28]
  PIN i2c_master.pwdata[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 12.7125 39.3900 12.7875 39.9000 ;
    END
  END i2c_master.pwdata[27]
  PIN i2c_master.pwdata[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 30.4125 0.5100 30.4875 ;
    END
  END i2c_master.pwdata[26]
  PIN i2c_master.pwdata[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 11.3625 39.3900 11.4375 39.9000 ;
    END
  END i2c_master.pwdata[25]
  PIN i2c_master.pwdata[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 28.9125 39.3900 28.9875 39.9000 ;
    END
  END i2c_master.pwdata[24]
  PIN i2c_master.pwdata[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 30.7125 0.5100 30.7875 ;
    END
  END i2c_master.pwdata[23]
  PIN i2c_master.pwdata[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10.4625 39.3900 10.5375 39.9000 ;
    END
  END i2c_master.pwdata[22]
  PIN i2c_master.pwdata[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 31.0125 0.5100 31.0875 ;
    END
  END i2c_master.pwdata[21]
  PIN i2c_master.pwdata[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 31.0125 0.5100 31.0875 ;
    END
  END i2c_master.pwdata[20]
  PIN i2c_master.pwdata[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 17.3625 0.0000 17.4375 0.5100 ;
    END
  END i2c_master.pwdata[19]
  PIN i2c_master.pwdata[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 36.4125 0.5100 36.4875 ;
    END
  END i2c_master.pwdata[18]
  PIN i2c_master.pwdata[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 10.0125 0.5100 10.0875 ;
    END
  END i2c_master.pwdata[17]
  PIN i2c_master.pwdata[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5.3175 39.4800 5.3925 39.9000 ;
    END
  END i2c_master.pwdata[16]
  PIN i2c_master.pwdata[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15.6075 0.0000 15.6825 0.4200 ;
    END
  END i2c_master.pwdata[15]
  PIN i2c_master.pwdata[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10.1625 0.0000 10.2375 0.5100 ;
    END
  END i2c_master.pwdata[14]
  PIN i2c_master.pwdata[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 14.2125 0.0000 14.2875 0.5100 ;
    END
  END i2c_master.pwdata[13]
  PIN i2c_master.pwdata[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 10.0125 0.5100 10.0875 ;
    END
  END i2c_master.pwdata[12]
  PIN i2c_master.pwdata[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11.0625 39.3900 11.1375 39.9000 ;
    END
  END i2c_master.pwdata[11]
  PIN i2c_master.pwdata[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 9.7125 0.5100 9.7875 ;
    END
  END i2c_master.pwdata[10]
  PIN i2c_master.pwdata[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 31.3125 0.5100 31.3875 ;
    END
  END i2c_master.pwdata[9]
  PIN i2c_master.pwdata[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 11.0625 39.3900 11.1375 39.9000 ;
    END
  END i2c_master.pwdata[8]
  PIN i2c_master.pwdata[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 9.7125 0.5100 9.7875 ;
    END
  END i2c_master.pwdata[7]
  PIN i2c_master.pwdata[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 13.6125 0.0000 13.6875 0.5100 ;
    END
  END i2c_master.pwdata[6]
  PIN i2c_master.pwdata[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 29.3625 39.3900 29.4375 39.9000 ;
    END
  END i2c_master.pwdata[5]
  PIN i2c_master.pwdata[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 0.0000 9.3000 2.1225 9.9000 ;
    END
  END i2c_master.pwdata[4]
  PIN i2c_master.pwdata[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 9.4125 0.5100 9.4875 ;
    END
  END i2c_master.pwdata[3]
  PIN i2c_master.pwdata[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 9.4125 0.5100 9.4875 ;
    END
  END i2c_master.pwdata[2]
  PIN i2c_master.pwdata[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 9.1125 0.5100 9.1875 ;
    END
  END i2c_master.pwdata[1]
  PIN i2c_master.pwdata[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10.7625 39.3900 10.8375 39.9000 ;
    END
  END i2c_master.pwdata[0]
  PIN i2c_master.pwrite
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4.6875 0.0000 4.7625 0.4200 ;
    END
  END i2c_master.pwrite
  PIN i2c_master.psel
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 21.4875 0.0000 21.5625 0.4200 ;
    END
  END i2c_master.psel
  PIN i2c_master.penable
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 2.8125 0.5100 2.8875 ;
    END
  END i2c_master.penable
  PIN i2c_master.prdata[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 20.9625 39.3900 21.0375 39.9000 ;
    END
  END i2c_master.prdata[31]
  PIN i2c_master.prdata[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 25.6125 39.3900 25.6875 39.9000 ;
    END
  END i2c_master.prdata[30]
  PIN i2c_master.prdata[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.8100 34.7625 40.3200 34.8375 ;
    END
  END i2c_master.prdata[29]
  PIN i2c_master.prdata[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.8100 8.5125 40.3200 8.5875 ;
    END
  END i2c_master.prdata[28]
  PIN i2c_master.prdata[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 38.1975 8.1000 40.3200 8.7000 ;
    END
  END i2c_master.prdata[27]
  PIN i2c_master.prdata[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 18.8625 39.3900 18.9375 39.9000 ;
    END
  END i2c_master.prdata[26]
  PIN i2c_master.prdata[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 27.4125 39.3900 27.4875 39.9000 ;
    END
  END i2c_master.prdata[25]
  PIN i2c_master.prdata[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 28.1625 39.3900 28.2375 39.9000 ;
    END
  END i2c_master.prdata[24]
  PIN i2c_master.prdata[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 30.5625 39.3900 30.6375 39.9000 ;
    END
  END i2c_master.prdata[23]
  PIN i2c_master.prdata[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.8100 35.0625 40.3200 35.1375 ;
    END
  END i2c_master.prdata[22]
  PIN i2c_master.prdata[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.8100 8.2125 40.3200 8.2875 ;
    END
  END i2c_master.prdata[21]
  PIN i2c_master.prdata[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.8100 35.3625 40.3200 35.4375 ;
    END
  END i2c_master.prdata[20]
  PIN i2c_master.prdata[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.8100 35.6625 40.3200 35.7375 ;
    END
  END i2c_master.prdata[19]
  PIN i2c_master.prdata[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.8100 7.9125 40.3200 7.9875 ;
    END
  END i2c_master.prdata[18]
  PIN i2c_master.prdata[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 28.3125 39.3900 28.3875 39.9000 ;
    END
  END i2c_master.prdata[17]
  PIN i2c_master.prdata[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 25.9125 39.3900 25.9875 39.9000 ;
    END
  END i2c_master.prdata[16]
  PIN i2c_master.prdata[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 26.2125 39.3900 26.2875 39.9000 ;
    END
  END i2c_master.prdata[15]
  PIN i2c_master.prdata[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 22.9125 39.3900 22.9875 39.9000 ;
    END
  END i2c_master.prdata[14]
  PIN i2c_master.prdata[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.8100 7.6125 40.3200 7.6875 ;
    END
  END i2c_master.prdata[13]
  PIN i2c_master.prdata[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 33.7125 39.3900 33.7875 39.9000 ;
    END
  END i2c_master.prdata[12]
  PIN i2c_master.prdata[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 26.8125 39.3900 26.8875 39.9000 ;
    END
  END i2c_master.prdata[11]
  PIN i2c_master.prdata[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 23.0625 39.3900 23.1375 39.9000 ;
    END
  END i2c_master.prdata[10]
  PIN i2c_master.prdata[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.8100 7.3125 40.3200 7.3875 ;
    END
  END i2c_master.prdata[9]
  PIN i2c_master.prdata[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 13.0125 39.3900 13.0875 39.9000 ;
    END
  END i2c_master.prdata[8]
  PIN i2c_master.prdata[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 37.2375 39.4800 37.3125 39.9000 ;
    END
  END i2c_master.prdata[7]
  PIN i2c_master.prdata[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.8100 35.9625 40.3200 36.0375 ;
    END
  END i2c_master.prdata[6]
  PIN i2c_master.prdata[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 23.6625 39.3900 23.7375 39.9000 ;
    END
  END i2c_master.prdata[5]
  PIN i2c_master.prdata[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 26.5125 39.3900 26.5875 39.9000 ;
    END
  END i2c_master.prdata[4]
  PIN i2c_master.prdata[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 35.7675 39.4800 35.8425 39.9000 ;
    END
  END i2c_master.prdata[3]
  PIN i2c_master.prdata[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 33.8775 39.4800 33.9525 39.9000 ;
    END
  END i2c_master.prdata[2]
  PIN i2c_master.prdata[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 29.2125 39.3900 29.2875 39.9000 ;
    END
  END i2c_master.prdata[1]
  PIN i2c_master.prdata[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.8100 7.0125 40.3200 7.0875 ;
    END
  END i2c_master.prdata[0]
  PIN i2c_master.pready
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 35.8125 0.0000 35.8875 0.5100 ;
    END
  END i2c_master.pready
  PIN i2c_master.pslverr
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 30.8625 0.0000 30.9375 0.5100 ;
    END
  END i2c_master.pslverr
  PIN fll_master.paddr[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 27.5625 40.3200 27.6375 ;
    END
  END fll_master.paddr[31]
  PIN fll_master.paddr[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 27.8625 40.3200 27.9375 ;
    END
  END fll_master.paddr[30]
  PIN fll_master.paddr[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 28.1625 40.3200 28.2375 ;
    END
  END fll_master.paddr[29]
  PIN fll_master.paddr[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16.9125 0.0000 16.9875 0.5100 ;
    END
  END fll_master.paddr[28]
  PIN fll_master.paddr[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17.2125 0.0000 17.2875 0.5100 ;
    END
  END fll_master.paddr[27]
  PIN fll_master.paddr[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 28.4625 40.3200 28.5375 ;
    END
  END fll_master.paddr[26]
  PIN fll_master.paddr[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17.5125 0.0000 17.5875 0.5100 ;
    END
  END fll_master.paddr[25]
  PIN fll_master.paddr[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 28.7625 40.3200 28.8375 ;
    END
  END fll_master.paddr[24]
  PIN fll_master.paddr[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 29.0625 40.3200 29.1375 ;
    END
  END fll_master.paddr[23]
  PIN fll_master.paddr[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 29.3625 40.3200 29.4375 ;
    END
  END fll_master.paddr[22]
  PIN fll_master.paddr[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 29.6625 40.3200 29.7375 ;
    END
  END fll_master.paddr[21]
  PIN fll_master.paddr[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17.8125 0.0000 17.8875 0.5100 ;
    END
  END fll_master.paddr[20]
  PIN fll_master.paddr[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 29.9625 40.3200 30.0375 ;
    END
  END fll_master.paddr[19]
  PIN fll_master.paddr[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 30.2625 40.3200 30.3375 ;
    END
  END fll_master.paddr[18]
  PIN fll_master.paddr[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 30.5625 40.3200 30.6375 ;
    END
  END fll_master.paddr[17]
  PIN fll_master.paddr[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 30.8625 40.3200 30.9375 ;
    END
  END fll_master.paddr[16]
  PIN fll_master.paddr[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 31.1625 40.3200 31.2375 ;
    END
  END fll_master.paddr[15]
  PIN fll_master.paddr[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18.1125 0.0000 18.1875 0.5100 ;
    END
  END fll_master.paddr[14]
  PIN fll_master.paddr[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18.4125 0.0000 18.4875 0.5100 ;
    END
  END fll_master.paddr[13]
  PIN fll_master.paddr[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 31.4625 40.3200 31.5375 ;
    END
  END fll_master.paddr[12]
  PIN fll_master.paddr[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8.0625 39.3900 8.1375 39.9000 ;
    END
  END fll_master.paddr[11]
  PIN fll_master.paddr[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 22.7625 0.5100 22.8375 ;
    END
  END fll_master.paddr[10]
  PIN fll_master.paddr[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8.8875 39.4800 8.9625 39.9000 ;
    END
  END fll_master.paddr[9]
  PIN fll_master.paddr[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13.7625 39.3900 13.8375 39.9000 ;
    END
  END fll_master.paddr[8]
  PIN fll_master.paddr[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 0.0000 26.1000 2.1225 26.7000 ;
    END
  END fll_master.paddr[7]
  PIN fll_master.paddr[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14.0625 39.3900 14.1375 39.9000 ;
    END
  END fll_master.paddr[6]
  PIN fll_master.paddr[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 23.0625 0.5100 23.1375 ;
    END
  END fll_master.paddr[5]
  PIN fll_master.paddr[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 13.9125 0.5100 13.9875 ;
    END
  END fll_master.paddr[4]
  PIN fll_master.paddr[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 29.8125 0.5100 29.8875 ;
    END
  END fll_master.paddr[3]
  PIN fll_master.paddr[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15.1125 39.3900 15.1875 39.9000 ;
    END
  END fll_master.paddr[2]
  PIN fll_master.paddr[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12.4575 39.4800 12.5325 39.9000 ;
    END
  END fll_master.paddr[1]
  PIN fll_master.paddr[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8.8125 39.3900 8.8875 39.9000 ;
    END
  END fll_master.paddr[0]
  PIN fll_master.pwdata[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 19.6125 0.5100 19.6875 ;
    END
  END fll_master.pwdata[31]
  PIN fll_master.pwdata[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 13.9125 0.5100 13.9875 ;
    END
  END fll_master.pwdata[30]
  PIN fll_master.pwdata[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 34.3125 0.5100 34.3875 ;
    END
  END fll_master.pwdata[29]
  PIN fll_master.pwdata[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 13.6125 0.5100 13.6875 ;
    END
  END fll_master.pwdata[28]
  PIN fll_master.pwdata[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 17.6625 39.3900 17.7375 39.9000 ;
    END
  END fll_master.pwdata[27]
  PIN fll_master.pwdata[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 30.7125 0.5100 30.7875 ;
    END
  END fll_master.pwdata[26]
  PIN fll_master.pwdata[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 11.9625 39.3900 12.0375 39.9000 ;
    END
  END fll_master.pwdata[25]
  PIN fll_master.pwdata[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 19.1625 39.3900 19.2375 39.9000 ;
    END
  END fll_master.pwdata[24]
  PIN fll_master.pwdata[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 21.4125 0.5100 21.4875 ;
    END
  END fll_master.pwdata[23]
  PIN fll_master.pwdata[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 26.8125 0.5100 26.8875 ;
    END
  END fll_master.pwdata[22]
  PIN fll_master.pwdata[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 24.4125 0.5100 24.4875 ;
    END
  END fll_master.pwdata[21]
  PIN fll_master.pwdata[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 21.2625 0.5100 21.3375 ;
    END
  END fll_master.pwdata[20]
  PIN fll_master.pwdata[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 19.3125 0.5100 19.3875 ;
    END
  END fll_master.pwdata[19]
  PIN fll_master.pwdata[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 34.0125 0.5100 34.0875 ;
    END
  END fll_master.pwdata[18]
  PIN fll_master.pwdata[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 20.8125 0.5100 20.8875 ;
    END
  END fll_master.pwdata[17]
  PIN fll_master.pwdata[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6.4125 39.3900 6.4875 39.9000 ;
    END
  END fll_master.pwdata[16]
  PIN fll_master.pwdata[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17.2125 39.3900 17.2875 39.9000 ;
    END
  END fll_master.pwdata[15]
  PIN fll_master.pwdata[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 19.0125 0.5100 19.0875 ;
    END
  END fll_master.pwdata[14]
  PIN fll_master.pwdata[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 16.6125 0.5100 16.6875 ;
    END
  END fll_master.pwdata[13]
  PIN fll_master.pwdata[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 21.1125 0.5100 21.1875 ;
    END
  END fll_master.pwdata[12]
  PIN fll_master.pwdata[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15.6075 39.4800 15.6825 39.9000 ;
    END
  END fll_master.pwdata[11]
  PIN fll_master.pwdata[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 14.2125 0.5100 14.2875 ;
    END
  END fll_master.pwdata[10]
  PIN fll_master.pwdata[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 28.3125 0.5100 28.3875 ;
    END
  END fll_master.pwdata[9]
  PIN fll_master.pwdata[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 16.1625 39.3900 16.2375 39.9000 ;
    END
  END fll_master.pwdata[8]
  PIN fll_master.pwdata[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 18.4125 0.5100 18.4875 ;
    END
  END fll_master.pwdata[7]
  PIN fll_master.pwdata[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 15.4125 0.5100 15.4875 ;
    END
  END fll_master.pwdata[6]
  PIN fll_master.pwdata[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18.4125 39.3900 18.4875 39.9000 ;
    END
  END fll_master.pwdata[5]
  PIN fll_master.pwdata[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 13.6125 0.5100 13.6875 ;
    END
  END fll_master.pwdata[4]
  PIN fll_master.pwdata[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 14.2125 0.5100 14.2875 ;
    END
  END fll_master.pwdata[3]
  PIN fll_master.pwdata[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 18.5625 0.5100 18.6375 ;
    END
  END fll_master.pwdata[2]
  PIN fll_master.pwdata[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 0.0000 14.1000 2.1225 14.7000 ;
    END
  END fll_master.pwdata[1]
  PIN fll_master.pwdata[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 26.2125 0.5100 26.2875 ;
    END
  END fll_master.pwdata[0]
  PIN fll_master.pwrite
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 2.5125 0.5100 2.5875 ;
    END
  END fll_master.pwrite
  PIN fll_master.psel
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18.3375 0.0000 18.4125 0.4200 ;
    END
  END fll_master.psel
  PIN fll_master.penable
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 2.5125 0.5100 2.5875 ;
    END
  END fll_master.penable
  PIN fll_master.prdata[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 22.1625 39.3900 22.2375 39.9000 ;
    END
  END fll_master.prdata[31]
  PIN fll_master.prdata[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 24.7125 39.3900 24.7875 39.9000 ;
    END
  END fll_master.prdata[30]
  PIN fll_master.prdata[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.8100 29.6625 40.3200 29.7375 ;
    END
  END fll_master.prdata[29]
  PIN fll_master.prdata[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.8100 18.2625 40.3200 18.3375 ;
    END
  END fll_master.prdata[28]
  PIN fll_master.prdata[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.8100 11.2125 40.3200 11.2875 ;
    END
  END fll_master.prdata[27]
  PIN fll_master.prdata[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 22.7625 39.3900 22.8375 39.9000 ;
    END
  END fll_master.prdata[26]
  PIN fll_master.prdata[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 27.1125 39.3900 27.1875 39.9000 ;
    END
  END fll_master.prdata[25]
  PIN fll_master.prdata[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 26.9475 39.4800 27.0225 39.9000 ;
    END
  END fll_master.prdata[24]
  PIN fll_master.prdata[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.8100 27.2625 40.3200 27.3375 ;
    END
  END fll_master.prdata[23]
  PIN fll_master.prdata[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.8100 29.3625 40.3200 29.4375 ;
    END
  END fll_master.prdata[22]
  PIN fll_master.prdata[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.8100 17.9625 40.3200 18.0375 ;
    END
  END fll_master.prdata[21]
  PIN fll_master.prdata[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.8100 30.2625 40.3200 30.3375 ;
    END
  END fll_master.prdata[20]
  PIN fll_master.prdata[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 38.1975 30.9000 40.3200 31.5000 ;
    END
  END fll_master.prdata[19]
  PIN fll_master.prdata[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.8100 20.9625 40.3200 21.0375 ;
    END
  END fll_master.prdata[18]
  PIN fll_master.prdata[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.8100 20.3625 40.3200 20.4375 ;
    END
  END fll_master.prdata[17]
  PIN fll_master.prdata[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 24.7125 39.3900 24.7875 39.9000 ;
    END
  END fll_master.prdata[16]
  PIN fll_master.prdata[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.8100 24.1125 40.3200 24.1875 ;
    END
  END fll_master.prdata[15]
  PIN fll_master.prdata[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.8100 10.9125 40.3200 10.9875 ;
    END
  END fll_master.prdata[14]
  PIN fll_master.prdata[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 38.1975 10.5000 40.3200 11.1000 ;
    END
  END fll_master.prdata[13]
  PIN fll_master.prdata[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 30.1125 39.3900 30.1875 39.9000 ;
    END
  END fll_master.prdata[12]
  PIN fll_master.prdata[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 29.6625 39.3900 29.7375 39.9000 ;
    END
  END fll_master.prdata[11]
  PIN fll_master.prdata[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 22.3125 39.3900 22.3875 39.9000 ;
    END
  END fll_master.prdata[10]
  PIN fll_master.prdata[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.8100 10.6125 40.3200 10.6875 ;
    END
  END fll_master.prdata[9]
  PIN fll_master.prdata[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 22.0125 39.3900 22.0875 39.9000 ;
    END
  END fll_master.prdata[8]
  PIN fll_master.prdata[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 32.3625 39.3900 32.4375 39.9000 ;
    END
  END fll_master.prdata[7]
  PIN fll_master.prdata[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.8100 31.4625 40.3200 31.5375 ;
    END
  END fll_master.prdata[6]
  PIN fll_master.prdata[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 22.4625 39.3900 22.5375 39.9000 ;
    END
  END fll_master.prdata[5]
  PIN fll_master.prdata[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 25.4775 39.4800 25.5525 39.9000 ;
    END
  END fll_master.prdata[4]
  PIN fll_master.prdata[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.8100 31.7625 40.3200 31.8375 ;
    END
  END fll_master.prdata[3]
  PIN fll_master.prdata[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 27.5625 39.3900 27.6375 39.9000 ;
    END
  END fll_master.prdata[2]
  PIN fll_master.prdata[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 29.2575 39.4800 29.3325 39.9000 ;
    END
  END fll_master.prdata[1]
  PIN fll_master.prdata[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.8100 10.3125 40.3200 10.3875 ;
    END
  END fll_master.prdata[0]
  PIN fll_master.pready
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 32.4075 0.0000 32.4825 0.4200 ;
    END
  END fll_master.pready
  PIN fll_master.pslverr
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 29.8875 0.0000 29.9625 0.4200 ;
    END
  END fll_master.pslverr
  PIN soc_ctrl_master.paddr[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 31.7625 40.3200 31.8375 ;
    END
  END soc_ctrl_master.paddr[31]
  PIN soc_ctrl_master.paddr[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 32.0625 40.3200 32.1375 ;
    END
  END soc_ctrl_master.paddr[30]
  PIN soc_ctrl_master.paddr[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 32.3625 40.3200 32.4375 ;
    END
  END soc_ctrl_master.paddr[29]
  PIN soc_ctrl_master.paddr[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.8100 11.8125 40.3200 11.8875 ;
    END
  END soc_ctrl_master.paddr[28]
  PIN soc_ctrl_master.paddr[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.8100 12.1125 40.3200 12.1875 ;
    END
  END soc_ctrl_master.paddr[27]
  PIN soc_ctrl_master.paddr[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 32.6625 40.3200 32.7375 ;
    END
  END soc_ctrl_master.paddr[26]
  PIN soc_ctrl_master.paddr[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.8100 12.4125 40.3200 12.4875 ;
    END
  END soc_ctrl_master.paddr[25]
  PIN soc_ctrl_master.paddr[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 32.9625 40.3200 33.0375 ;
    END
  END soc_ctrl_master.paddr[24]
  PIN soc_ctrl_master.paddr[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 33.2625 40.3200 33.3375 ;
    END
  END soc_ctrl_master.paddr[23]
  PIN soc_ctrl_master.paddr[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 33.5625 40.3200 33.6375 ;
    END
  END soc_ctrl_master.paddr[22]
  PIN soc_ctrl_master.paddr[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 33.8625 40.3200 33.9375 ;
    END
  END soc_ctrl_master.paddr[21]
  PIN soc_ctrl_master.paddr[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.8100 12.7125 40.3200 12.7875 ;
    END
  END soc_ctrl_master.paddr[20]
  PIN soc_ctrl_master.paddr[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 34.1625 40.3200 34.2375 ;
    END
  END soc_ctrl_master.paddr[19]
  PIN soc_ctrl_master.paddr[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 34.4625 40.3200 34.5375 ;
    END
  END soc_ctrl_master.paddr[18]
  PIN soc_ctrl_master.paddr[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 34.7625 40.3200 34.8375 ;
    END
  END soc_ctrl_master.paddr[17]
  PIN soc_ctrl_master.paddr[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 35.0625 40.3200 35.1375 ;
    END
  END soc_ctrl_master.paddr[16]
  PIN soc_ctrl_master.paddr[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 35.3625 40.3200 35.4375 ;
    END
  END soc_ctrl_master.paddr[15]
  PIN soc_ctrl_master.paddr[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.8100 13.0125 40.3200 13.0875 ;
    END
  END soc_ctrl_master.paddr[14]
  PIN soc_ctrl_master.paddr[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.8100 13.3125 40.3200 13.3875 ;
    END
  END soc_ctrl_master.paddr[13]
  PIN soc_ctrl_master.paddr[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.8100 13.6125 40.3200 13.6875 ;
    END
  END soc_ctrl_master.paddr[12]
  PIN soc_ctrl_master.paddr[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7.6275 39.4800 7.7025 39.9000 ;
    END
  END soc_ctrl_master.paddr[11]
  PIN soc_ctrl_master.paddr[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 31.3125 0.5100 31.3875 ;
    END
  END soc_ctrl_master.paddr[10]
  PIN soc_ctrl_master.paddr[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8.5125 39.3900 8.5875 39.9000 ;
    END
  END soc_ctrl_master.paddr[9]
  PIN soc_ctrl_master.paddr[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 10.7625 39.3900 10.8375 39.9000 ;
    END
  END soc_ctrl_master.paddr[8]
  PIN soc_ctrl_master.paddr[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 31.6125 0.5100 31.6875 ;
    END
  END soc_ctrl_master.paddr[7]
  PIN soc_ctrl_master.paddr[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 9.2625 39.3900 9.3375 39.9000 ;
    END
  END soc_ctrl_master.paddr[6]
  PIN soc_ctrl_master.paddr[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 8.9625 39.3900 9.0375 39.9000 ;
    END
  END soc_ctrl_master.paddr[5]
  PIN soc_ctrl_master.paddr[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 9.1125 0.5100 9.1875 ;
    END
  END soc_ctrl_master.paddr[4]
  PIN soc_ctrl_master.paddr[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 31.6125 0.5100 31.6875 ;
    END
  END soc_ctrl_master.paddr[3]
  PIN soc_ctrl_master.paddr[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 8.6625 39.3900 8.7375 39.9000 ;
    END
  END soc_ctrl_master.paddr[2]
  PIN soc_ctrl_master.paddr[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 7.9125 39.3900 7.9875 39.9000 ;
    END
  END soc_ctrl_master.paddr[1]
  PIN soc_ctrl_master.paddr[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 7.6125 39.3900 7.6875 39.9000 ;
    END
  END soc_ctrl_master.paddr[0]
  PIN soc_ctrl_master.pwdata[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 12.4125 0.0000 12.4875 0.5100 ;
    END
  END soc_ctrl_master.pwdata[31]
  PIN soc_ctrl_master.pwdata[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10.9125 0.0000 10.9875 0.5100 ;
    END
  END soc_ctrl_master.pwdata[30]
  PIN soc_ctrl_master.pwdata[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 32.2125 0.5100 32.2875 ;
    END
  END soc_ctrl_master.pwdata[29]
  PIN soc_ctrl_master.pwdata[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 8.8125 0.5100 8.8875 ;
    END
  END soc_ctrl_master.pwdata[28]
  PIN soc_ctrl_master.pwdata[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7.4625 39.3900 7.5375 39.9000 ;
    END
  END soc_ctrl_master.pwdata[27]
  PIN soc_ctrl_master.pwdata[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 0.0000 32.1000 2.1225 32.7000 ;
    END
  END soc_ctrl_master.pwdata[26]
  PIN soc_ctrl_master.pwdata[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 32.5125 0.5100 32.5875 ;
    END
  END soc_ctrl_master.pwdata[25]
  PIN soc_ctrl_master.pwdata[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 32.5125 39.3900 32.5875 39.9000 ;
    END
  END soc_ctrl_master.pwdata[24]
  PIN soc_ctrl_master.pwdata[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 33.1125 0.5100 33.1875 ;
    END
  END soc_ctrl_master.pwdata[23]
  PIN soc_ctrl_master.pwdata[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 7.3125 39.3900 7.3875 39.9000 ;
    END
  END soc_ctrl_master.pwdata[22]
  PIN soc_ctrl_master.pwdata[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 33.4125 0.5100 33.4875 ;
    END
  END soc_ctrl_master.pwdata[21]
  PIN soc_ctrl_master.pwdata[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 33.4125 0.5100 33.4875 ;
    END
  END soc_ctrl_master.pwdata[20]
  PIN soc_ctrl_master.pwdata[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 19.1625 0.0000 19.2375 0.5100 ;
    END
  END soc_ctrl_master.pwdata[19]
  PIN soc_ctrl_master.pwdata[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4.0125 39.3900 4.0875 39.9000 ;
    END
  END soc_ctrl_master.pwdata[18]
  PIN soc_ctrl_master.pwdata[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 8.8125 0.5100 8.8875 ;
    END
  END soc_ctrl_master.pwdata[17]
  PIN soc_ctrl_master.pwdata[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5.9475 39.4800 6.0225 39.9000 ;
    END
  END soc_ctrl_master.pwdata[16]
  PIN soc_ctrl_master.pwdata[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16.6575 0.0000 16.7325 0.4200 ;
    END
  END soc_ctrl_master.pwdata[15]
  PIN soc_ctrl_master.pwdata[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11.6175 0.0000 11.6925 0.4200 ;
    END
  END soc_ctrl_master.pwdata[14]
  PIN soc_ctrl_master.pwdata[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12.7125 0.0000 12.7875 0.5100 ;
    END
  END soc_ctrl_master.pwdata[13]
  PIN soc_ctrl_master.pwdata[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 8.5125 0.5100 8.5875 ;
    END
  END soc_ctrl_master.pwdata[12]
  PIN soc_ctrl_master.pwdata[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13.4625 0.0000 13.5375 0.5100 ;
    END
  END soc_ctrl_master.pwdata[11]
  PIN soc_ctrl_master.pwdata[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 8.5125 0.5100 8.5875 ;
    END
  END soc_ctrl_master.pwdata[10]
  PIN soc_ctrl_master.pwdata[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 33.7125 0.5100 33.7875 ;
    END
  END soc_ctrl_master.pwdata[9]
  PIN soc_ctrl_master.pwdata[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 7.0125 39.3900 7.0875 39.9000 ;
    END
  END soc_ctrl_master.pwdata[8]
  PIN soc_ctrl_master.pwdata[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8.8125 0.0000 8.8875 0.5100 ;
    END
  END soc_ctrl_master.pwdata[7]
  PIN soc_ctrl_master.pwdata[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 12.8625 0.0000 12.9375 0.5100 ;
    END
  END soc_ctrl_master.pwdata[6]
  PIN soc_ctrl_master.pwdata[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 19.7625 0.0000 19.8375 0.5100 ;
    END
  END soc_ctrl_master.pwdata[5]
  PIN soc_ctrl_master.pwdata[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9.3075 0.0000 9.3825 0.4200 ;
    END
  END soc_ctrl_master.pwdata[4]
  PIN soc_ctrl_master.pwdata[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 8.2125 0.5100 8.2875 ;
    END
  END soc_ctrl_master.pwdata[3]
  PIN soc_ctrl_master.pwdata[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 8.2125 0.5100 8.2875 ;
    END
  END soc_ctrl_master.pwdata[2]
  PIN soc_ctrl_master.pwdata[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 7.9125 0.5100 7.9875 ;
    END
  END soc_ctrl_master.pwdata[1]
  PIN soc_ctrl_master.pwdata[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6.7875 39.4800 6.8625 39.9000 ;
    END
  END soc_ctrl_master.pwdata[0]
  PIN soc_ctrl_master.pwrite
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 2.2125 0.5100 2.2875 ;
    END
  END soc_ctrl_master.pwrite
  PIN soc_ctrl_master.psel
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.8100 13.9125 40.3200 13.9875 ;
    END
  END soc_ctrl_master.psel
  PIN soc_ctrl_master.penable
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 2.2125 0.5100 2.2875 ;
    END
  END soc_ctrl_master.penable
  PIN soc_ctrl_master.prdata[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 29.9625 39.3900 30.0375 39.9000 ;
    END
  END soc_ctrl_master.prdata[31]
  PIN soc_ctrl_master.prdata[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 30.7275 39.4800 30.8025 39.9000 ;
    END
  END soc_ctrl_master.prdata[30]
  PIN soc_ctrl_master.prdata[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 36.6075 39.4800 36.6825 39.9000 ;
    END
  END soc_ctrl_master.prdata[29]
  PIN soc_ctrl_master.prdata[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.8100 6.7125 40.3200 6.7875 ;
    END
  END soc_ctrl_master.prdata[28]
  PIN soc_ctrl_master.prdata[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.8100 6.4125 40.3200 6.4875 ;
    END
  END soc_ctrl_master.prdata[27]
  PIN soc_ctrl_master.prdata[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 30.2625 39.3900 30.3375 39.9000 ;
    END
  END soc_ctrl_master.prdata[26]
  PIN soc_ctrl_master.prdata[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 30.5625 39.3900 30.6375 39.9000 ;
    END
  END soc_ctrl_master.prdata[25]
  PIN soc_ctrl_master.prdata[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 30.8625 39.3900 30.9375 39.9000 ;
    END
  END soc_ctrl_master.prdata[24]
  PIN soc_ctrl_master.prdata[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 31.1625 39.3900 31.2375 39.9000 ;
    END
  END soc_ctrl_master.prdata[23]
  PIN soc_ctrl_master.prdata[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.8100 36.2625 40.3200 36.3375 ;
    END
  END soc_ctrl_master.prdata[22]
  PIN soc_ctrl_master.prdata[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.8100 6.1125 40.3200 6.1875 ;
    END
  END soc_ctrl_master.prdata[21]
  PIN soc_ctrl_master.prdata[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 36.4125 39.3900 36.4875 39.9000 ;
    END
  END soc_ctrl_master.prdata[20]
  PIN soc_ctrl_master.prdata[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 36.1125 39.3900 36.1875 39.9000 ;
    END
  END soc_ctrl_master.prdata[19]
  PIN soc_ctrl_master.prdata[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.8100 36.5625 40.3200 36.6375 ;
    END
  END soc_ctrl_master.prdata[18]
  PIN soc_ctrl_master.prdata[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 30.8625 39.3900 30.9375 39.9000 ;
    END
  END soc_ctrl_master.prdata[17]
  PIN soc_ctrl_master.prdata[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 31.4625 39.3900 31.5375 39.9000 ;
    END
  END soc_ctrl_master.prdata[16]
  PIN soc_ctrl_master.prdata[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 22.5375 0.0000 22.6125 0.4200 ;
    END
  END soc_ctrl_master.prdata[15]
  PIN soc_ctrl_master.prdata[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 21.1125 0.0000 21.1875 0.5100 ;
    END
  END soc_ctrl_master.prdata[14]
  PIN soc_ctrl_master.prdata[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.8100 5.5125 40.3200 5.5875 ;
    END
  END soc_ctrl_master.prdata[13]
  PIN soc_ctrl_master.prdata[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 32.6625 39.3900 32.7375 39.9000 ;
    END
  END soc_ctrl_master.prdata[12]
  PIN soc_ctrl_master.prdata[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 31.6125 39.3900 31.6875 39.9000 ;
    END
  END soc_ctrl_master.prdata[11]
  PIN soc_ctrl_master.prdata[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 31.9125 0.5100 31.9875 ;
    END
  END soc_ctrl_master.prdata[10]
  PIN soc_ctrl_master.prdata[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.8100 5.2125 40.3200 5.2875 ;
    END
  END soc_ctrl_master.prdata[9]
  PIN soc_ctrl_master.prdata[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 31.9125 0.5100 31.9875 ;
    END
  END soc_ctrl_master.prdata[8]
  PIN soc_ctrl_master.prdata[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 35.8125 39.3900 35.8875 39.9000 ;
    END
  END soc_ctrl_master.prdata[7]
  PIN soc_ctrl_master.prdata[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.8100 36.8625 40.3200 36.9375 ;
    END
  END soc_ctrl_master.prdata[6]
  PIN soc_ctrl_master.prdata[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 31.1625 39.3900 31.2375 39.9000 ;
    END
  END soc_ctrl_master.prdata[5]
  PIN soc_ctrl_master.prdata[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 31.9125 39.3900 31.9875 39.9000 ;
    END
  END soc_ctrl_master.prdata[4]
  PIN soc_ctrl_master.prdata[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.8100 37.6125 40.3200 37.6875 ;
    END
  END soc_ctrl_master.prdata[3]
  PIN soc_ctrl_master.prdata[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 34.2975 39.4800 34.3725 39.9000 ;
    END
  END soc_ctrl_master.prdata[2]
  PIN soc_ctrl_master.prdata[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 32.2125 39.3900 32.2875 39.9000 ;
    END
  END soc_ctrl_master.prdata[1]
  PIN soc_ctrl_master.prdata[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.8100 4.9125 40.3200 4.9875 ;
    END
  END soc_ctrl_master.prdata[0]
  PIN soc_ctrl_master.pready
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 36.8625 0.0000 36.9375 0.5100 ;
    END
  END soc_ctrl_master.pready
  PIN soc_ctrl_master.pslverr
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 28.9125 0.0000 28.9875 0.5100 ;
    END
  END soc_ctrl_master.pslverr
  PIN debug_master.paddr[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 35.6625 40.3200 35.7375 ;
    END
  END debug_master.paddr[31]
  PIN debug_master.paddr[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 35.9625 40.3200 36.0375 ;
    END
  END debug_master.paddr[30]
  PIN debug_master.paddr[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 36.2625 40.3200 36.3375 ;
    END
  END debug_master.paddr[29]
  PIN debug_master.paddr[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 23.5125 0.0000 23.5875 0.5100 ;
    END
  END debug_master.paddr[28]
  PIN debug_master.paddr[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 23.8125 0.0000 23.8875 0.5100 ;
    END
  END debug_master.paddr[27]
  PIN debug_master.paddr[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 36.5625 40.3200 36.6375 ;
    END
  END debug_master.paddr[26]
  PIN debug_master.paddr[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 24.1125 0.0000 24.1875 0.5100 ;
    END
  END debug_master.paddr[25]
  PIN debug_master.paddr[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 36.8625 40.3200 36.9375 ;
    END
  END debug_master.paddr[24]
  PIN debug_master.paddr[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 37.1625 40.3200 37.2375 ;
    END
  END debug_master.paddr[23]
  PIN debug_master.paddr[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 37.4625 40.3200 37.5375 ;
    END
  END debug_master.paddr[22]
  PIN debug_master.paddr[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 37.7625 40.3200 37.8375 ;
    END
  END debug_master.paddr[21]
  PIN debug_master.paddr[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 24.4125 0.0000 24.4875 0.5100 ;
    END
  END debug_master.paddr[20]
  PIN debug_master.paddr[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 38.0625 40.3200 38.1375 ;
    END
  END debug_master.paddr[19]
  PIN debug_master.paddr[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 38.3625 40.3200 38.4375 ;
    END
  END debug_master.paddr[18]
  PIN debug_master.paddr[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 38.6625 40.3200 38.7375 ;
    END
  END debug_master.paddr[17]
  PIN debug_master.paddr[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 24.7125 0.0000 24.7875 0.5100 ;
    END
  END debug_master.paddr[16]
  PIN debug_master.paddr[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.8100 38.9625 40.3200 39.0375 ;
    END
  END debug_master.paddr[15]
  PIN debug_master.paddr[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 25.0125 0.0000 25.0875 0.5100 ;
    END
  END debug_master.paddr[14]
  PIN debug_master.paddr[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 26.3175 0.0000 26.3925 0.4200 ;
    END
  END debug_master.paddr[13]
  PIN debug_master.paddr[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 25.3125 0.0000 25.3875 0.5100 ;
    END
  END debug_master.paddr[12]
  PIN debug_master.paddr[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7.2075 39.4800 7.2825 39.9000 ;
    END
  END debug_master.paddr[11]
  PIN debug_master.paddr[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 23.8125 0.5100 23.8875 ;
    END
  END debug_master.paddr[10]
  PIN debug_master.paddr[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10.1625 39.3900 10.2375 39.9000 ;
    END
  END debug_master.paddr[9]
  PIN debug_master.paddr[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14.5125 39.3900 14.5875 39.9000 ;
    END
  END debug_master.paddr[8]
  PIN debug_master.paddr[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 28.0125 0.5100 28.0875 ;
    END
  END debug_master.paddr[7]
  PIN debug_master.paddr[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13.5075 39.4800 13.5825 39.9000 ;
    END
  END debug_master.paddr[6]
  PIN debug_master.paddr[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 23.8125 0.5100 23.8875 ;
    END
  END debug_master.paddr[5]
  PIN debug_master.paddr[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 11.8125 0.5100 11.8875 ;
    END
  END debug_master.paddr[4]
  PIN debug_master.paddr[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 28.6125 0.5100 28.6875 ;
    END
  END debug_master.paddr[3]
  PIN debug_master.paddr[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15.1875 39.4800 15.2625 39.9000 ;
    END
  END debug_master.paddr[2]
  PIN debug_master.paddr[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11.9625 39.3900 12.0375 39.9000 ;
    END
  END debug_master.paddr[1]
  PIN debug_master.paddr[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9.7125 39.3900 9.7875 39.9000 ;
    END
  END debug_master.paddr[0]
  PIN debug_master.pwdata[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 19.6125 0.5100 19.6875 ;
    END
  END debug_master.pwdata[31]
  PIN debug_master.pwdata[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 11.8125 0.5100 11.8875 ;
    END
  END debug_master.pwdata[30]
  PIN debug_master.pwdata[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 32.8125 0.5100 32.8875 ;
    END
  END debug_master.pwdata[29]
  PIN debug_master.pwdata[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 0.0000 11.7000 2.1225 12.3000 ;
    END
  END debug_master.pwdata[28]
  PIN debug_master.pwdata[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18.1125 39.3900 18.1875 39.9000 ;
    END
  END debug_master.pwdata[27]
  PIN debug_master.pwdata[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 30.1125 0.5100 30.1875 ;
    END
  END debug_master.pwdata[26]
  PIN debug_master.pwdata[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 12.2625 39.3900 12.3375 39.9000 ;
    END
  END debug_master.pwdata[25]
  PIN debug_master.pwdata[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 19.7625 39.3900 19.8375 39.9000 ;
    END
  END debug_master.pwdata[24]
  PIN debug_master.pwdata[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 0.0000 23.7000 2.1225 24.3000 ;
    END
  END debug_master.pwdata[23]
  PIN debug_master.pwdata[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 28.0125 0.5100 28.0875 ;
    END
  END debug_master.pwdata[22]
  PIN debug_master.pwdata[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 25.9125 0.5100 25.9875 ;
    END
  END debug_master.pwdata[21]
  PIN debug_master.pwdata[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 21.7125 0.5100 21.7875 ;
    END
  END debug_master.pwdata[20]
  PIN debug_master.pwdata[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 20.2125 0.5100 20.2875 ;
    END
  END debug_master.pwdata[19]
  PIN debug_master.pwdata[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 34.9125 0.5100 34.9875 ;
    END
  END debug_master.pwdata[18]
  PIN debug_master.pwdata[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 0.0000 20.1000 2.1225 20.7000 ;
    END
  END debug_master.pwdata[17]
  PIN debug_master.pwdata[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6.1125 39.3900 6.1875 39.9000 ;
    END
  END debug_master.pwdata[16]
  PIN debug_master.pwdata[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17.7075 39.4800 17.7825 39.9000 ;
    END
  END debug_master.pwdata[15]
  PIN debug_master.pwdata[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 18.1125 0.5100 18.1875 ;
    END
  END debug_master.pwdata[14]
  PIN debug_master.pwdata[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 17.5125 0.5100 17.5875 ;
    END
  END debug_master.pwdata[13]
  PIN debug_master.pwdata[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 22.1625 0.5100 22.2375 ;
    END
  END debug_master.pwdata[12]
  PIN debug_master.pwdata[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 21.5625 0.5100 21.6375 ;
    END
  END debug_master.pwdata[11]
  PIN debug_master.pwdata[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 11.2125 0.5100 11.2875 ;
    END
  END debug_master.pwdata[10]
  PIN debug_master.pwdata[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 26.5125 0.5100 26.5875 ;
    END
  END debug_master.pwdata[9]
  PIN debug_master.pwdata[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15.4125 39.3900 15.4875 39.9000 ;
    END
  END debug_master.pwdata[8]
  PIN debug_master.pwdata[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 17.3625 0.5100 17.4375 ;
    END
  END debug_master.pwdata[7]
  PIN debug_master.pwdata[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14.1375 0.0000 14.2125 0.4200 ;
    END
  END debug_master.pwdata[6]
  PIN debug_master.pwdata[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18.9675 39.4800 19.0425 39.9000 ;
    END
  END debug_master.pwdata[5]
  PIN debug_master.pwdata[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 11.5125 0.5100 11.5875 ;
    END
  END debug_master.pwdata[4]
  PIN debug_master.pwdata[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 11.5125 0.5100 11.5875 ;
    END
  END debug_master.pwdata[3]
  PIN debug_master.pwdata[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 17.2125 0.5100 17.2875 ;
    END
  END debug_master.pwdata[2]
  PIN debug_master.pwdata[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 11.2125 0.5100 11.2875 ;
    END
  END debug_master.pwdata[1]
  PIN debug_master.pwdata[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11.6175 39.4800 11.6925 39.9000 ;
    END
  END debug_master.pwdata[0]
  PIN debug_master.pwrite
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2.7975 0.0000 2.8725 0.4200 ;
    END
  END debug_master.pwrite
  PIN debug_master.psel
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 24.6375 0.0000 24.7125 0.4200 ;
    END
  END debug_master.psel
  PIN debug_master.penable
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1.9125 0.5100 1.9875 ;
    END
  END debug_master.penable
  PIN debug_master.prdata[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 23.7975 39.4800 23.8725 39.9000 ;
    END
  END debug_master.prdata[31]
  PIN debug_master.prdata[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 25.0575 39.4800 25.1325 39.9000 ;
    END
  END debug_master.prdata[30]
  PIN debug_master.prdata[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.8100 28.7625 40.3200 28.8375 ;
    END
  END debug_master.prdata[29]
  PIN debug_master.prdata[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.8100 19.4625 40.3200 19.5375 ;
    END
  END debug_master.prdata[28]
  PIN debug_master.prdata[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.8100 15.2625 40.3200 15.3375 ;
    END
  END debug_master.prdata[27]
  PIN debug_master.prdata[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 23.1675 39.4800 23.2425 39.9000 ;
    END
  END debug_master.prdata[26]
  PIN debug_master.prdata[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 27.3675 39.4800 27.4425 39.9000 ;
    END
  END debug_master.prdata[25]
  PIN debug_master.prdata[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 26.3175 39.4800 26.3925 39.9000 ;
    END
  END debug_master.prdata[24]
  PIN debug_master.prdata[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 28.4175 39.4800 28.4925 39.9000 ;
    END
  END debug_master.prdata[23]
  PIN debug_master.prdata[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.8100 28.0125 40.3200 28.0875 ;
    END
  END debug_master.prdata[22]
  PIN debug_master.prdata[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.8100 17.3625 40.3200 17.4375 ;
    END
  END debug_master.prdata[21]
  PIN debug_master.prdata[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.8100 28.3125 40.3200 28.3875 ;
    END
  END debug_master.prdata[20]
  PIN debug_master.prdata[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.8100 30.8625 40.3200 30.9375 ;
    END
  END debug_master.prdata[19]
  PIN debug_master.prdata[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.8100 23.5125 40.3200 23.5875 ;
    END
  END debug_master.prdata[18]
  PIN debug_master.prdata[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.8100 16.7625 40.3200 16.8375 ;
    END
  END debug_master.prdata[17]
  PIN debug_master.prdata[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 25.0125 39.3900 25.0875 39.9000 ;
    END
  END debug_master.prdata[16]
  PIN debug_master.prdata[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.8100 16.1625 40.3200 16.2375 ;
    END
  END debug_master.prdata[15]
  PIN debug_master.prdata[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.8100 16.4625 40.3200 16.5375 ;
    END
  END debug_master.prdata[14]
  PIN debug_master.prdata[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.8100 14.2125 40.3200 14.2875 ;
    END
  END debug_master.prdata[13]
  PIN debug_master.prdata[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.8100 30.5625 40.3200 30.6375 ;
    END
  END debug_master.prdata[12]
  PIN debug_master.prdata[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.8100 24.4125 40.3200 24.4875 ;
    END
  END debug_master.prdata[11]
  PIN debug_master.prdata[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 23.9625 39.3900 24.0375 39.9000 ;
    END
  END debug_master.prdata[10]
  PIN debug_master.prdata[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.8100 21.5625 40.3200 21.6375 ;
    END
  END debug_master.prdata[9]
  PIN debug_master.prdata[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 24.4125 39.3900 24.4875 39.9000 ;
    END
  END debug_master.prdata[8]
  PIN debug_master.prdata[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 31.7775 39.4800 31.8525 39.9000 ;
    END
  END debug_master.prdata[7]
  PIN debug_master.prdata[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.8100 23.2125 40.3200 23.2875 ;
    END
  END debug_master.prdata[6]
  PIN debug_master.prdata[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 23.3625 39.3900 23.4375 39.9000 ;
    END
  END debug_master.prdata[5]
  PIN debug_master.prdata[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 26.3625 39.3900 26.4375 39.9000 ;
    END
  END debug_master.prdata[4]
  PIN debug_master.prdata[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.8100 26.0625 40.3200 26.1375 ;
    END
  END debug_master.prdata[3]
  PIN debug_master.prdata[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 28.0125 39.3900 28.0875 39.9000 ;
    END
  END debug_master.prdata[2]
  PIN debug_master.prdata[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 28.8375 39.4800 28.9125 39.9000 ;
    END
  END debug_master.prdata[1]
  PIN debug_master.prdata[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.8100 15.8625 40.3200 15.9375 ;
    END
  END debug_master.prdata[0]
  PIN debug_master.pready
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 31.5675 0.0000 31.6425 0.4200 ;
    END
  END debug_master.pready
  PIN debug_master.pslverr
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 30.1125 0.0000 30.1875 0.5100 ;
    END
  END debug_master.pslverr
  OBS
    LAYER M1 ;
        RECT 0.0000 0.0000 40.3200 39.9000 ;
    LAYER M2 ;
        RECT 0.0000 0.0000 40.3200 39.9000 ;
    LAYER M3 ;
        RECT 0.0000 0.0000 40.3200 39.9000 ;
    LAYER M4 ;
        RECT 0.0000 0.0000 40.3200 39.9000 ;
    LAYER M5 ;
        RECT 0.0000 0.0000 40.3200 39.9000 ;
    LAYER M6 ;
        RECT 0.0000 0.0000 40.3200 39.9000 ;
    LAYER M7 ;
        RECT 0.0000 0.0000 40.3200 39.9000 ;
    LAYER M8 ;
        RECT 0.0000 0.0000 40.3200 39.9000 ;
  END
END periph_bus_wrap


